module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module add(clk, add_a, add_b, add_z);
  input clk;
  input [31:0] add_a;
  input [31:0] add_b;
  output [31:0] add_z;
  wire [31:0] s_0;
  wire [31:0] s_1;
  wire [31:0] s_2;
  wire [0:0] s_3;
  wire [0:0] s_4;
  wire [0:0] s_5;
  wire [0:0] s_6;
  wire [0:0] s_7;
  wire [0:0] s_8;
  wire [31:0] s_9;
  wire [0:0] s_10;
  wire [31:0] s_11;
  wire [0:0] s_12;
  wire [0:0] s_13;
  wire [0:0] s_14;
  wire [8:0] s_15;
  wire [7:0] s_16;
  wire [7:0] s_17;
  wire [7:0] s_18;
  wire [7:0] s_19;
  wire [6:0] s_20;
  wire [0:0] s_21;
  wire [7:0] s_22;
  wire [8:0] s_23;
  wire [7:0] s_24;
  wire [7:0] s_25;
  wire [7:0] s_26;
  wire [7:0] s_27;
  wire [6:0] s_28;
  wire [0:0] s_29;
  wire [7:0] s_30;
  wire [0:0] s_31;
  wire [0:0] s_32;
  wire [7:0] s_33;
  wire [0:0] s_34;
  wire [22:0] s_35;
  wire [22:0] s_36;
  wire [0:0] s_37;
  wire [0:0] s_38;
  wire [0:0] s_39;
  wire [7:0] s_40;
  wire [0:0] s_41;
  wire [22:0] s_42;
  wire [22:0] s_43;
  wire [0:0] s_44;
  wire [0:0] s_45;
  wire [27:0] s_46;
  wire [27:0] s_47;
  wire [23:0] s_48;
  wire [23:0] s_49;
  wire [0:0] s_50;
  wire [0:0] s_51;
  wire [0:0] s_52;
  wire [23:0] s_53;
  wire [0:0] s_54;
  wire [0:0] s_55;
  wire [0:0] s_56;
  wire [1:0] s_57;
  wire [27:0] s_58;
  wire [27:0] s_59;
  wire [27:0] s_60;
  wire [27:0] s_61;
  wire [23:0] s_62;
  wire [1:0] s_63;
  wire [8:0] s_64;
  wire [8:0] s_65;
  wire [8:0] s_66;
  wire [0:0] s_67;
  wire [27:0] s_68;
  wire [27:0] s_69;
  wire [27:0] s_70;
  wire [0:0] s_71;
  wire [0:0] s_72;
  wire [27:0] s_73;
  wire [27:0] s_74;
  wire [27:0] s_75;
  wire [27:0] s_76;
  wire [27:0] s_77;
  wire [27:0] s_78;
  wire [27:0] s_79;
  wire [27:0] s_80;
  wire [27:0] s_81;
  wire [0:0] s_82;
  wire [0:0] s_83;
  wire [30:0] s_84;
  wire [31:0] s_85;
  wire [31:0] s_86;
  wire [31:0] s_87;
  wire [30:0] s_88;
  wire [31:0] s_89;
  wire [31:0] s_90;
  wire [31:0] s_91;
  wire [30:0] s_92;
  wire [31:0] s_93;
  wire [31:0] s_94;
  wire [8:0] s_95;
  wire [8:0] s_96;
  wire [7:0] s_97;
  wire [22:0] s_98;
  wire [23:0] s_99;
  wire [23:0] s_100;
  wire [23:0] s_101;
  wire [24:0] s_102;
  wire [24:0] s_103;
  wire [24:0] s_104;
  wire [24:0] s_105;
  wire [23:0] s_106;
  wire [27:0] s_107;
  wire [27:0] s_108;
  wire [27:0] s_109;
  wire [27:0] s_110;
  wire [8:0] s_111;
  wire [8:0] s_112;
  wire [5:0] s_113;
  wire [5:0] s_114;
  wire [0:0] s_115;
  wire [0:0] s_116;
  wire [4:0] s_117;
  wire [0:0] s_118;
  wire [0:0] s_119;
  wire [3:0] s_120;
  wire [0:0] s_121;
  wire [0:0] s_122;
  wire [2:0] s_123;
  wire [0:0] s_124;
  wire [0:0] s_125;
  wire [1:0] s_126;
  wire [0:0] s_127;
  wire [0:0] s_128;
  wire [0:0] s_129;
  wire [1:0] s_130;
  wire [3:0] s_131;
  wire [7:0] s_132;
  wire [15:0] s_133;
  wire [31:0] s_134;
  wire [30:0] s_135;
  wire [29:0] s_136;
  wire [28:0] s_137;
  wire [0:0] s_138;
  wire [0:0] s_139;
  wire [0:0] s_140;
  wire [0:0] s_141;
  wire [0:0] s_142;
  wire [0:0] s_143;
  wire [0:0] s_144;
  wire [0:0] s_145;
  wire [0:0] s_146;
  wire [0:0] s_147;
  wire [0:0] s_148;
  wire [1:0] s_149;
  wire [0:0] s_150;
  wire [0:0] s_151;
  wire [0:0] s_152;
  wire [1:0] s_153;
  wire [0:0] s_154;
  wire [0:0] s_155;
  wire [0:0] s_156;
  wire [0:0] s_157;
  wire [0:0] s_158;
  wire [0:0] s_159;
  wire [1:0] s_160;
  wire [0:0] s_161;
  wire [0:0] s_162;
  wire [0:0] s_163;
  wire [0:0] s_164;
  wire [0:0] s_165;
  wire [0:0] s_166;
  wire [2:0] s_167;
  wire [0:0] s_168;
  wire [0:0] s_169;
  wire [1:0] s_170;
  wire [0:0] s_171;
  wire [0:0] s_172;
  wire [0:0] s_173;
  wire [1:0] s_174;
  wire [3:0] s_175;
  wire [0:0] s_176;
  wire [0:0] s_177;
  wire [0:0] s_178;
  wire [0:0] s_179;
  wire [0:0] s_180;
  wire [0:0] s_181;
  wire [0:0] s_182;
  wire [1:0] s_183;
  wire [0:0] s_184;
  wire [0:0] s_185;
  wire [0:0] s_186;
  wire [1:0] s_187;
  wire [0:0] s_188;
  wire [0:0] s_189;
  wire [0:0] s_190;
  wire [0:0] s_191;
  wire [0:0] s_192;
  wire [0:0] s_193;
  wire [1:0] s_194;
  wire [0:0] s_195;
  wire [0:0] s_196;
  wire [0:0] s_197;
  wire [0:0] s_198;
  wire [0:0] s_199;
  wire [2:0] s_200;
  wire [0:0] s_201;
  wire [0:0] s_202;
  wire [1:0] s_203;
  wire [1:0] s_204;
  wire [1:0] s_205;
  wire [0:0] s_206;
  wire [3:0] s_207;
  wire [0:0] s_208;
  wire [0:0] s_209;
  wire [2:0] s_210;
  wire [0:0] s_211;
  wire [0:0] s_212;
  wire [1:0] s_213;
  wire [0:0] s_214;
  wire [0:0] s_215;
  wire [0:0] s_216;
  wire [1:0] s_217;
  wire [3:0] s_218;
  wire [7:0] s_219;
  wire [0:0] s_220;
  wire [0:0] s_221;
  wire [0:0] s_222;
  wire [0:0] s_223;
  wire [0:0] s_224;
  wire [0:0] s_225;
  wire [0:0] s_226;
  wire [1:0] s_227;
  wire [0:0] s_228;
  wire [0:0] s_229;
  wire [0:0] s_230;
  wire [1:0] s_231;
  wire [0:0] s_232;
  wire [0:0] s_233;
  wire [0:0] s_234;
  wire [0:0] s_235;
  wire [0:0] s_236;
  wire [0:0] s_237;
  wire [1:0] s_238;
  wire [0:0] s_239;
  wire [0:0] s_240;
  wire [0:0] s_241;
  wire [0:0] s_242;
  wire [0:0] s_243;
  wire [0:0] s_244;
  wire [2:0] s_245;
  wire [0:0] s_246;
  wire [0:0] s_247;
  wire [1:0] s_248;
  wire [0:0] s_249;
  wire [0:0] s_250;
  wire [0:0] s_251;
  wire [1:0] s_252;
  wire [3:0] s_253;
  wire [0:0] s_254;
  wire [0:0] s_255;
  wire [0:0] s_256;
  wire [0:0] s_257;
  wire [0:0] s_258;
  wire [0:0] s_259;
  wire [0:0] s_260;
  wire [1:0] s_261;
  wire [0:0] s_262;
  wire [0:0] s_263;
  wire [0:0] s_264;
  wire [1:0] s_265;
  wire [0:0] s_266;
  wire [0:0] s_267;
  wire [0:0] s_268;
  wire [0:0] s_269;
  wire [0:0] s_270;
  wire [0:0] s_271;
  wire [1:0] s_272;
  wire [0:0] s_273;
  wire [0:0] s_274;
  wire [0:0] s_275;
  wire [0:0] s_276;
  wire [0:0] s_277;
  wire [2:0] s_278;
  wire [0:0] s_279;
  wire [0:0] s_280;
  wire [1:0] s_281;
  wire [1:0] s_282;
  wire [1:0] s_283;
  wire [3:0] s_284;
  wire [0:0] s_285;
  wire [0:0] s_286;
  wire [2:0] s_287;
  wire [2:0] s_288;
  wire [2:0] s_289;
  wire [0:0] s_290;
  wire [4:0] s_291;
  wire [0:0] s_292;
  wire [0:0] s_293;
  wire [3:0] s_294;
  wire [0:0] s_295;
  wire [0:0] s_296;
  wire [2:0] s_297;
  wire [0:0] s_298;
  wire [0:0] s_299;
  wire [1:0] s_300;
  wire [0:0] s_301;
  wire [0:0] s_302;
  wire [0:0] s_303;
  wire [1:0] s_304;
  wire [3:0] s_305;
  wire [7:0] s_306;
  wire [15:0] s_307;
  wire [0:0] s_308;
  wire [0:0] s_309;
  wire [0:0] s_310;
  wire [0:0] s_311;
  wire [0:0] s_312;
  wire [0:0] s_313;
  wire [0:0] s_314;
  wire [1:0] s_315;
  wire [0:0] s_316;
  wire [0:0] s_317;
  wire [0:0] s_318;
  wire [1:0] s_319;
  wire [0:0] s_320;
  wire [0:0] s_321;
  wire [0:0] s_322;
  wire [0:0] s_323;
  wire [0:0] s_324;
  wire [0:0] s_325;
  wire [1:0] s_326;
  wire [0:0] s_327;
  wire [0:0] s_328;
  wire [0:0] s_329;
  wire [0:0] s_330;
  wire [0:0] s_331;
  wire [0:0] s_332;
  wire [2:0] s_333;
  wire [0:0] s_334;
  wire [0:0] s_335;
  wire [1:0] s_336;
  wire [0:0] s_337;
  wire [0:0] s_338;
  wire [0:0] s_339;
  wire [1:0] s_340;
  wire [3:0] s_341;
  wire [0:0] s_342;
  wire [0:0] s_343;
  wire [0:0] s_344;
  wire [0:0] s_345;
  wire [0:0] s_346;
  wire [0:0] s_347;
  wire [0:0] s_348;
  wire [1:0] s_349;
  wire [0:0] s_350;
  wire [0:0] s_351;
  wire [0:0] s_352;
  wire [1:0] s_353;
  wire [0:0] s_354;
  wire [0:0] s_355;
  wire [0:0] s_356;
  wire [0:0] s_357;
  wire [0:0] s_358;
  wire [0:0] s_359;
  wire [1:0] s_360;
  wire [0:0] s_361;
  wire [0:0] s_362;
  wire [0:0] s_363;
  wire [0:0] s_364;
  wire [0:0] s_365;
  wire [2:0] s_366;
  wire [0:0] s_367;
  wire [0:0] s_368;
  wire [1:0] s_369;
  wire [1:0] s_370;
  wire [1:0] s_371;
  wire [0:0] s_372;
  wire [3:0] s_373;
  wire [0:0] s_374;
  wire [0:0] s_375;
  wire [2:0] s_376;
  wire [0:0] s_377;
  wire [0:0] s_378;
  wire [1:0] s_379;
  wire [0:0] s_380;
  wire [0:0] s_381;
  wire [0:0] s_382;
  wire [1:0] s_383;
  wire [3:0] s_384;
  wire [7:0] s_385;
  wire [0:0] s_386;
  wire [0:0] s_387;
  wire [0:0] s_388;
  wire [0:0] s_389;
  wire [0:0] s_390;
  wire [0:0] s_391;
  wire [0:0] s_392;
  wire [1:0] s_393;
  wire [0:0] s_394;
  wire [0:0] s_395;
  wire [0:0] s_396;
  wire [1:0] s_397;
  wire [0:0] s_398;
  wire [0:0] s_399;
  wire [0:0] s_400;
  wire [0:0] s_401;
  wire [0:0] s_402;
  wire [0:0] s_403;
  wire [1:0] s_404;
  wire [0:0] s_405;
  wire [0:0] s_406;
  wire [0:0] s_407;
  wire [0:0] s_408;
  wire [0:0] s_409;
  wire [0:0] s_410;
  wire [2:0] s_411;
  wire [0:0] s_412;
  wire [0:0] s_413;
  wire [1:0] s_414;
  wire [0:0] s_415;
  wire [0:0] s_416;
  wire [0:0] s_417;
  wire [1:0] s_418;
  wire [3:0] s_419;
  wire [0:0] s_420;
  wire [0:0] s_421;
  wire [0:0] s_422;
  wire [0:0] s_423;
  wire [0:0] s_424;
  wire [0:0] s_425;
  wire [0:0] s_426;
  wire [1:0] s_427;
  wire [0:0] s_428;
  wire [0:0] s_429;
  wire [0:0] s_430;
  wire [1:0] s_431;
  wire [0:0] s_432;
  wire [0:0] s_433;
  wire [0:0] s_434;
  wire [0:0] s_435;
  wire [0:0] s_436;
  wire [0:0] s_437;
  wire [1:0] s_438;
  wire [0:0] s_439;
  wire [0:0] s_440;
  wire [0:0] s_441;
  wire [0:0] s_442;
  wire [0:0] s_443;
  wire [2:0] s_444;
  wire [0:0] s_445;
  wire [0:0] s_446;
  wire [1:0] s_447;
  wire [1:0] s_448;
  wire [1:0] s_449;
  wire [3:0] s_450;
  wire [0:0] s_451;
  wire [0:0] s_452;
  wire [2:0] s_453;
  wire [2:0] s_454;
  wire [2:0] s_455;
  wire [4:0] s_456;
  wire [0:0] s_457;
  wire [0:0] s_458;
  wire [3:0] s_459;
  wire [3:0] s_460;
  wire [3:0] s_461;
  wire [8:0] s_462;
  wire [8:0] s_463;
  wire [8:0] s_464;
  wire [8:0] s_465;
  wire [8:0] s_466;
  wire [8:0] s_467;
  wire [0:0] s_468;
  wire [8:0] s_469;
  wire [0:0] s_470;
  wire [8:0] s_471;
  wire [8:0] s_472;
  wire [0:0] s_473;
  wire [23:0] s_474;
  wire [0:0] s_475;
  wire [0:0] s_476;
  wire [0:0] s_477;
  wire [0:0] s_478;
  wire [0:0] s_479;
  wire [0:0] s_480;
  wire [0:0] s_481;
  wire [0:0] s_482;
  wire [0:0] s_483;
  wire [0:0] s_484;
  wire [0:0] s_485;
  wire [0:0] s_486;
  wire [0:0] s_487;
  wire [23:0] s_488;
  wire [0:0] s_489;
  wire [31:0] s_490;
  wire [8:0] s_491;
  wire [0:0] s_492;
  wire [7:0] s_493;
  wire [7:0] s_494;
  wire [8:0] s_495;
  wire [8:0] s_496;
  wire [8:0] s_497;
  wire [8:0] s_498;
  wire [8:0] s_499;
  wire [8:0] s_500;
  wire [6:0] s_501;
  wire [22:0] s_502;
  wire [0:0] s_503;
  wire [0:0] s_504;
  wire [7:0] s_505;
  wire [0:0] s_506;
  wire [0:0] s_507;
  wire [0:0] s_508;
  wire [23:0] s_509;
  wire [0:0] s_510;
  wire [0:0] s_511;
  wire [0:0] s_512;
  wire [7:0] s_513;
  wire [0:0] s_514;
  wire [0:0] s_515;
  wire [0:0] s_516;
  wire [0:0] s_517;
  wire [0:0] s_518;
  wire [0:0] s_519;
  wire [0:0] s_520;
  wire [7:0] s_521;
  wire [0:0] s_522;
  wire [22:0] s_523;
  wire [0:0] s_524;
  wire [0:0] s_525;
  wire [7:0] s_526;
  wire [0:0] s_527;
  wire [22:0] s_528;
  wire [0:0] s_529;

  assign s_0 = s_516?s_1:s_85;
  dq #(32, 5) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_84};
  assign s_3 = s_72?s_4:s_5;
  assign s_4 = 1'd0;
  dq #(1, 2) dq_s_5 (clk, s_5, s_6);
  assign s_6 = s_45?s_7:s_44;
  assign s_7 = s_12?s_8:s_10;
  assign s_8 = s_9[31];
  assign s_9 = add_a;
  assign s_10 = s_11[31];
  assign s_11 = add_b;
  assign s_12 = s_13 & s_37;
  assign s_13 = s_14 | s_31;
  assign s_14 = $signed(s_15) > $signed(s_23);
  assign s_15 = $signed(s_16);
  assign s_16 = s_21?s_17:s_18;
  assign s_17 = -8'd126;
  assign s_18 = s_19 - s_20;
  assign s_19 = s_9[30:23];
  assign s_20 = 7'd127;
  assign s_21 = s_18 == s_22;
  assign s_22 = -8'd127;
  assign s_23 = $signed(s_24);
  assign s_24 = s_29?s_25:s_26;
  assign s_25 = -8'd126;
  assign s_26 = s_27 - s_28;
  assign s_27 = s_11[30:23];
  assign s_28 = 7'd127;
  assign s_29 = s_26 == s_30;
  assign s_30 = -8'd127;
  assign s_31 = s_32 & s_34;
  assign s_32 = s_18 == s_33;
  assign s_33 = 8'd128;
  assign s_34 = s_35 == s_36;
  assign s_35 = s_9[22:0];
  assign s_36 = 23'd0;
  assign s_37 = ~s_38;
  assign s_38 = s_39 & s_41;
  assign s_39 = s_26 == s_40;
  assign s_40 = 8'd128;
  assign s_41 = s_42 == s_43;
  assign s_42 = s_11[22:0];
  assign s_43 = 23'd0;
  assign s_44 = s_12?s_10:s_8;
  assign s_45 = s_46 >= s_58;
  assign s_46 = s_47 << s_57;
  assign s_47 = s_48;
  assign s_48 = s_12?s_49:s_53;
  assign s_49 = {s_50,s_35};
  assign s_50 = s_21?s_51:s_52;
  assign s_51 = 1'd0;
  assign s_52 = 1'd1;
  assign s_53 = {s_54,s_42};
  assign s_54 = s_29?s_55:s_56;
  assign s_55 = 1'd0;
  assign s_56 = 1'd1;
  assign s_57 = 2'd3;
  assign s_58 = s_59 | s_67;
  assign s_59 = s_60 >> s_64;
  assign s_60 = s_61 << s_63;
  assign s_61 = s_62;
  assign s_62 = s_12?s_53:s_49;
  assign s_63 = 2'd3;
  assign s_64 = s_65 - s_66;
  assign s_65 = s_12?s_15:s_23;
  assign s_66 = s_12?s_23:s_15;
  assign s_67 = s_68 != s_71;
  assign s_68 = s_60 << s_69;
  assign s_69 = s_70 - s_64;
  assign s_70 = 28'd28;
  assign s_71 = 1'd0;
  assign s_72 = s_73 == s_83;
  dq #(28, 1) dq_s_73 (clk, s_73, s_74);
  assign s_74 = s_75 + s_77;
  dq #(28, 1) dq_s_75 (clk, s_75, s_76);
  assign s_76 = s_45?s_46:s_58;
  dq #(28, 1) dq_s_77 (clk, s_77, s_78);
  assign s_78 = s_82?s_79:s_80;
  assign s_79 = s_45?s_58:s_46;
  assign s_80 = s_81 - s_79;
  assign s_81 = 28'd0;
  assign s_82 = s_8 == s_10;
  assign s_83 = 1'd0;
  assign s_84 = 31'd2143289344;
  assign s_85 = s_510?s_86:s_89;
  dq #(32, 5) dq_s_86 (clk, s_86, s_87);
  assign s_87 = {s_3,s_88};
  assign s_88 = 31'd2139095040;
  assign s_89 = s_508?s_90:s_93;
  dq #(32, 5) dq_s_90 (clk, s_90, s_91);
  assign s_91 = {s_3,s_92};
  assign s_92 = 31'd0;
  assign s_93 = s_503?s_94:s_490;
  assign s_94 = {s_95,s_98};
  dq #(9, 5) dq_s_95 (clk, s_95, s_96);
  assign s_96 = {s_3,s_97};
  assign s_97 = 8'd0;
  assign s_98 = s_99[22:0];
  dq #(24, 1) dq_s_99 (clk, s_99, s_100);
  assign s_100 = s_489?s_101:s_488;
  assign s_101 = s_102[24:1];
  assign s_102 = s_475?s_103:s_474;
  dq #(25, 1) dq_s_103 (clk, s_103, s_104);
  assign s_104 = s_105 + s_473;
  assign s_105 = s_106;
  assign s_106 = s_107[27:4];
  dq #(28, 1) dq_s_107 (clk, s_107, s_108);
  assign s_108 = s_109 << s_111;
  dq #(28, 2) dq_s_109 (clk, s_109, s_110);
  dq #(28, 1) dq_s_110 (clk, s_110, s_74);
  dq #(9, 1) dq_s_111 (clk, s_111, s_112);
  assign s_112 = s_470?s_113:s_462;
  dq #(6, 1) dq_s_113 (clk, s_113, s_114);
  assign s_114 = {s_115,s_456};
  assign s_115 = s_116 & s_290;
  assign s_116 = s_117[4];
  assign s_117 = {s_118,s_284};
  assign s_118 = s_119 & s_206;
  assign s_119 = s_120[3];
  assign s_120 = {s_121,s_200};
  assign s_121 = s_122 & s_166;
  assign s_122 = s_123[2];
  assign s_123 = {s_124,s_160};
  assign s_124 = s_125 & s_148;
  assign s_125 = s_126[1];
  assign s_126 = {s_127,s_144};
  assign s_127 = s_128 & s_142;
  assign s_128 = ~s_129;
  assign s_129 = s_130[1];
  assign s_130 = s_131[3:2];
  assign s_131 = s_132[7:4];
  assign s_132 = s_133[15:8];
  assign s_133 = s_134[31:16];
  assign s_134 = {s_135,s_141};
  assign s_135 = {s_136,s_140};
  assign s_136 = {s_137,s_139};
  assign s_137 = {s_110,s_138};
  assign s_138 = 1'd1;
  assign s_139 = 1'd1;
  assign s_140 = 1'd1;
  assign s_141 = 1'd1;
  assign s_142 = ~s_143;
  assign s_143 = s_130[0];
  assign s_144 = s_145 & s_147;
  assign s_145 = ~s_146;
  assign s_146 = s_130[1];
  assign s_147 = s_130[0];
  assign s_148 = s_149[1];
  assign s_149 = {s_150,s_156};
  assign s_150 = s_151 & s_154;
  assign s_151 = ~s_152;
  assign s_152 = s_153[1];
  assign s_153 = s_131[1:0];
  assign s_154 = ~s_155;
  assign s_155 = s_153[0];
  assign s_156 = s_157 & s_159;
  assign s_157 = ~s_158;
  assign s_158 = s_153[1];
  assign s_159 = s_153[0];
  assign s_160 = {s_161,s_163};
  assign s_161 = s_125 & s_162;
  assign s_162 = ~s_148;
  assign s_163 = s_125?s_164:s_165;
  assign s_164 = s_149[0:0];
  assign s_165 = s_126[0:0];
  assign s_166 = s_167[2];
  assign s_167 = {s_168,s_194};
  assign s_168 = s_169 & s_182;
  assign s_169 = s_170[1];
  assign s_170 = {s_171,s_178};
  assign s_171 = s_172 & s_176;
  assign s_172 = ~s_173;
  assign s_173 = s_174[1];
  assign s_174 = s_175[3:2];
  assign s_175 = s_132[3:0];
  assign s_176 = ~s_177;
  assign s_177 = s_174[0];
  assign s_178 = s_179 & s_181;
  assign s_179 = ~s_180;
  assign s_180 = s_174[1];
  assign s_181 = s_174[0];
  assign s_182 = s_183[1];
  assign s_183 = {s_184,s_190};
  assign s_184 = s_185 & s_188;
  assign s_185 = ~s_186;
  assign s_186 = s_187[1];
  assign s_187 = s_175[1:0];
  assign s_188 = ~s_189;
  assign s_189 = s_187[0];
  assign s_190 = s_191 & s_193;
  assign s_191 = ~s_192;
  assign s_192 = s_187[1];
  assign s_193 = s_187[0];
  assign s_194 = {s_195,s_197};
  assign s_195 = s_169 & s_196;
  assign s_196 = ~s_182;
  assign s_197 = s_169?s_198:s_199;
  assign s_198 = s_183[0:0];
  assign s_199 = s_170[0:0];
  assign s_200 = {s_201,s_203};
  assign s_201 = s_122 & s_202;
  assign s_202 = ~s_166;
  assign s_203 = s_122?s_204:s_205;
  assign s_204 = s_167[1:0];
  assign s_205 = s_123[1:0];
  assign s_206 = s_207[3];
  assign s_207 = {s_208,s_278};
  assign s_208 = s_209 & s_244;
  assign s_209 = s_210[2];
  assign s_210 = {s_211,s_238};
  assign s_211 = s_212 & s_226;
  assign s_212 = s_213[1];
  assign s_213 = {s_214,s_222};
  assign s_214 = s_215 & s_220;
  assign s_215 = ~s_216;
  assign s_216 = s_217[1];
  assign s_217 = s_218[3:2];
  assign s_218 = s_219[7:4];
  assign s_219 = s_133[7:0];
  assign s_220 = ~s_221;
  assign s_221 = s_217[0];
  assign s_222 = s_223 & s_225;
  assign s_223 = ~s_224;
  assign s_224 = s_217[1];
  assign s_225 = s_217[0];
  assign s_226 = s_227[1];
  assign s_227 = {s_228,s_234};
  assign s_228 = s_229 & s_232;
  assign s_229 = ~s_230;
  assign s_230 = s_231[1];
  assign s_231 = s_218[1:0];
  assign s_232 = ~s_233;
  assign s_233 = s_231[0];
  assign s_234 = s_235 & s_237;
  assign s_235 = ~s_236;
  assign s_236 = s_231[1];
  assign s_237 = s_231[0];
  assign s_238 = {s_239,s_241};
  assign s_239 = s_212 & s_240;
  assign s_240 = ~s_226;
  assign s_241 = s_212?s_242:s_243;
  assign s_242 = s_227[0:0];
  assign s_243 = s_213[0:0];
  assign s_244 = s_245[2];
  assign s_245 = {s_246,s_272};
  assign s_246 = s_247 & s_260;
  assign s_247 = s_248[1];
  assign s_248 = {s_249,s_256};
  assign s_249 = s_250 & s_254;
  assign s_250 = ~s_251;
  assign s_251 = s_252[1];
  assign s_252 = s_253[3:2];
  assign s_253 = s_219[3:0];
  assign s_254 = ~s_255;
  assign s_255 = s_252[0];
  assign s_256 = s_257 & s_259;
  assign s_257 = ~s_258;
  assign s_258 = s_252[1];
  assign s_259 = s_252[0];
  assign s_260 = s_261[1];
  assign s_261 = {s_262,s_268};
  assign s_262 = s_263 & s_266;
  assign s_263 = ~s_264;
  assign s_264 = s_265[1];
  assign s_265 = s_253[1:0];
  assign s_266 = ~s_267;
  assign s_267 = s_265[0];
  assign s_268 = s_269 & s_271;
  assign s_269 = ~s_270;
  assign s_270 = s_265[1];
  assign s_271 = s_265[0];
  assign s_272 = {s_273,s_275};
  assign s_273 = s_247 & s_274;
  assign s_274 = ~s_260;
  assign s_275 = s_247?s_276:s_277;
  assign s_276 = s_261[0:0];
  assign s_277 = s_248[0:0];
  assign s_278 = {s_279,s_281};
  assign s_279 = s_209 & s_280;
  assign s_280 = ~s_244;
  assign s_281 = s_209?s_282:s_283;
  assign s_282 = s_245[1:0];
  assign s_283 = s_210[1:0];
  assign s_284 = {s_285,s_287};
  assign s_285 = s_119 & s_286;
  assign s_286 = ~s_206;
  assign s_287 = s_119?s_288:s_289;
  assign s_288 = s_207[2:0];
  assign s_289 = s_120[2:0];
  assign s_290 = s_291[4];
  assign s_291 = {s_292,s_450};
  assign s_292 = s_293 & s_372;
  assign s_293 = s_294[3];
  assign s_294 = {s_295,s_366};
  assign s_295 = s_296 & s_332;
  assign s_296 = s_297[2];
  assign s_297 = {s_298,s_326};
  assign s_298 = s_299 & s_314;
  assign s_299 = s_300[1];
  assign s_300 = {s_301,s_310};
  assign s_301 = s_302 & s_308;
  assign s_302 = ~s_303;
  assign s_303 = s_304[1];
  assign s_304 = s_305[3:2];
  assign s_305 = s_306[7:4];
  assign s_306 = s_307[15:8];
  assign s_307 = s_134[15:0];
  assign s_308 = ~s_309;
  assign s_309 = s_304[0];
  assign s_310 = s_311 & s_313;
  assign s_311 = ~s_312;
  assign s_312 = s_304[1];
  assign s_313 = s_304[0];
  assign s_314 = s_315[1];
  assign s_315 = {s_316,s_322};
  assign s_316 = s_317 & s_320;
  assign s_317 = ~s_318;
  assign s_318 = s_319[1];
  assign s_319 = s_305[1:0];
  assign s_320 = ~s_321;
  assign s_321 = s_319[0];
  assign s_322 = s_323 & s_325;
  assign s_323 = ~s_324;
  assign s_324 = s_319[1];
  assign s_325 = s_319[0];
  assign s_326 = {s_327,s_329};
  assign s_327 = s_299 & s_328;
  assign s_328 = ~s_314;
  assign s_329 = s_299?s_330:s_331;
  assign s_330 = s_315[0:0];
  assign s_331 = s_300[0:0];
  assign s_332 = s_333[2];
  assign s_333 = {s_334,s_360};
  assign s_334 = s_335 & s_348;
  assign s_335 = s_336[1];
  assign s_336 = {s_337,s_344};
  assign s_337 = s_338 & s_342;
  assign s_338 = ~s_339;
  assign s_339 = s_340[1];
  assign s_340 = s_341[3:2];
  assign s_341 = s_306[3:0];
  assign s_342 = ~s_343;
  assign s_343 = s_340[0];
  assign s_344 = s_345 & s_347;
  assign s_345 = ~s_346;
  assign s_346 = s_340[1];
  assign s_347 = s_340[0];
  assign s_348 = s_349[1];
  assign s_349 = {s_350,s_356};
  assign s_350 = s_351 & s_354;
  assign s_351 = ~s_352;
  assign s_352 = s_353[1];
  assign s_353 = s_341[1:0];
  assign s_354 = ~s_355;
  assign s_355 = s_353[0];
  assign s_356 = s_357 & s_359;
  assign s_357 = ~s_358;
  assign s_358 = s_353[1];
  assign s_359 = s_353[0];
  assign s_360 = {s_361,s_363};
  assign s_361 = s_335 & s_362;
  assign s_362 = ~s_348;
  assign s_363 = s_335?s_364:s_365;
  assign s_364 = s_349[0:0];
  assign s_365 = s_336[0:0];
  assign s_366 = {s_367,s_369};
  assign s_367 = s_296 & s_368;
  assign s_368 = ~s_332;
  assign s_369 = s_296?s_370:s_371;
  assign s_370 = s_333[1:0];
  assign s_371 = s_297[1:0];
  assign s_372 = s_373[3];
  assign s_373 = {s_374,s_444};
  assign s_374 = s_375 & s_410;
  assign s_375 = s_376[2];
  assign s_376 = {s_377,s_404};
  assign s_377 = s_378 & s_392;
  assign s_378 = s_379[1];
  assign s_379 = {s_380,s_388};
  assign s_380 = s_381 & s_386;
  assign s_381 = ~s_382;
  assign s_382 = s_383[1];
  assign s_383 = s_384[3:2];
  assign s_384 = s_385[7:4];
  assign s_385 = s_307[7:0];
  assign s_386 = ~s_387;
  assign s_387 = s_383[0];
  assign s_388 = s_389 & s_391;
  assign s_389 = ~s_390;
  assign s_390 = s_383[1];
  assign s_391 = s_383[0];
  assign s_392 = s_393[1];
  assign s_393 = {s_394,s_400};
  assign s_394 = s_395 & s_398;
  assign s_395 = ~s_396;
  assign s_396 = s_397[1];
  assign s_397 = s_384[1:0];
  assign s_398 = ~s_399;
  assign s_399 = s_397[0];
  assign s_400 = s_401 & s_403;
  assign s_401 = ~s_402;
  assign s_402 = s_397[1];
  assign s_403 = s_397[0];
  assign s_404 = {s_405,s_407};
  assign s_405 = s_378 & s_406;
  assign s_406 = ~s_392;
  assign s_407 = s_378?s_408:s_409;
  assign s_408 = s_393[0:0];
  assign s_409 = s_379[0:0];
  assign s_410 = s_411[2];
  assign s_411 = {s_412,s_438};
  assign s_412 = s_413 & s_426;
  assign s_413 = s_414[1];
  assign s_414 = {s_415,s_422};
  assign s_415 = s_416 & s_420;
  assign s_416 = ~s_417;
  assign s_417 = s_418[1];
  assign s_418 = s_419[3:2];
  assign s_419 = s_385[3:0];
  assign s_420 = ~s_421;
  assign s_421 = s_418[0];
  assign s_422 = s_423 & s_425;
  assign s_423 = ~s_424;
  assign s_424 = s_418[1];
  assign s_425 = s_418[0];
  assign s_426 = s_427[1];
  assign s_427 = {s_428,s_434};
  assign s_428 = s_429 & s_432;
  assign s_429 = ~s_430;
  assign s_430 = s_431[1];
  assign s_431 = s_419[1:0];
  assign s_432 = ~s_433;
  assign s_433 = s_431[0];
  assign s_434 = s_435 & s_437;
  assign s_435 = ~s_436;
  assign s_436 = s_431[1];
  assign s_437 = s_431[0];
  assign s_438 = {s_439,s_441};
  assign s_439 = s_413 & s_440;
  assign s_440 = ~s_426;
  assign s_441 = s_413?s_442:s_443;
  assign s_442 = s_427[0:0];
  assign s_443 = s_414[0:0];
  assign s_444 = {s_445,s_447};
  assign s_445 = s_375 & s_446;
  assign s_446 = ~s_410;
  assign s_447 = s_375?s_448:s_449;
  assign s_448 = s_411[1:0];
  assign s_449 = s_376[1:0];
  assign s_450 = {s_451,s_453};
  assign s_451 = s_293 & s_452;
  assign s_452 = ~s_372;
  assign s_453 = s_293?s_454:s_455;
  assign s_454 = s_373[2:0];
  assign s_455 = s_294[2:0];
  assign s_456 = {s_457,s_459};
  assign s_457 = s_116 & s_458;
  assign s_458 = ~s_290;
  assign s_459 = s_116?s_460:s_461;
  assign s_460 = s_291[3:0];
  assign s_461 = s_117[3:0];
  dq #(9, 2) dq_s_462 (clk, s_462, s_463);
  assign s_463 = s_464 - s_469;
  dq #(9, 1) dq_s_464 (clk, s_464, s_465);
  assign s_465 = s_466 + s_468;
  assign s_466 = s_45?s_65:s_467;
  assign s_467 = s_66 + s_64;
  assign s_468 = 1'd1;
  assign s_469 = -9'd126;
  assign s_470 = s_471 <= s_472;
  assign s_471 = s_113;
  dq #(9, 2) dq_s_472 (clk, s_472, s_463);
  assign s_473 = 1'd1;
  dq #(24, 1) dq_s_474 (clk, s_474, s_106);
  assign s_475 = s_476 & s_478;
  dq #(1, 1) dq_s_476 (clk, s_476, s_477);
  assign s_477 = s_107[3];
  assign s_478 = s_479 | s_486;
  assign s_479 = s_480 | s_482;
  dq #(1, 1) dq_s_480 (clk, s_480, s_481);
  assign s_481 = s_107[2];
  dq #(1, 1) dq_s_482 (clk, s_482, s_483);
  assign s_483 = s_484 | s_485;
  assign s_484 = s_107[1];
  assign s_485 = s_107[0];
  dq #(1, 1) dq_s_486 (clk, s_486, s_487);
  assign s_487 = s_106[0];
  assign s_488 = s_102[23:0];
  assign s_489 = s_102[24];
  assign s_490 = {s_491,s_502};
  assign s_491 = {s_492,s_493};
  dq #(1, 5) dq_s_492 (clk, s_492, s_3);
  assign s_493 = s_494 + s_501;
  assign s_494 = s_495[7:0];
  dq #(9, 1) dq_s_495 (clk, s_495, s_496);
  assign s_496 = s_497 + s_489;
  dq #(9, 1) dq_s_497 (clk, s_497, s_498);
  dq #(9, 1) dq_s_498 (clk, s_498, s_499);
  assign s_499 = s_500 - s_111;
  dq #(9, 3) dq_s_500 (clk, s_500, s_464);
  assign s_501 = 7'd127;
  assign s_502 = s_99[22:0];
  assign s_503 = s_504 & s_506;
  assign s_504 = s_494 == s_505;
  assign s_505 = -8'd126;
  assign s_506 = ~s_507;
  assign s_507 = s_99[23];
  assign s_508 = s_99 == s_509;
  assign s_509 = 24'd0;
  assign s_510 = s_511 | s_515;
  assign s_511 = s_512 | s_514;
  assign s_512 = $signed(s_495) > $signed(s_513);
  assign s_513 = 8'd127;
  dq #(1, 7) dq_s_514 (clk, s_514, s_31);
  dq #(1, 7) dq_s_515 (clk, s_515, s_38);
  dq #(1, 7) dq_s_516 (clk, s_516, s_517);
  assign s_517 = s_518 | s_529;
  assign s_518 = s_519 | s_524;
  assign s_519 = s_520 & s_522;
  assign s_520 = s_18 == s_521;
  assign s_521 = 8'd128;
  assign s_522 = s_35 != s_523;
  assign s_523 = 23'd0;
  assign s_524 = s_525 & s_527;
  assign s_525 = s_26 == s_526;
  assign s_526 = 8'd128;
  assign s_527 = s_42 != s_528;
  assign s_528 = 23'd0;
  assign s_529 = s_31 & s_38;
  assign add_z = s_0;
endmodule
