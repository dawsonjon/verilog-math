module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module div(clk, div_a, div_b, div_z);
  input clk;
  input [31:0] div_a;
  input [31:0] div_b;
  output [31:0] div_z;
  wire [31:0] s_0;
  wire [31:0] s_1;
  wire [31:0] s_2;
  wire [0:0] s_3;
  wire [0:0] s_4;
  wire [31:0] s_5;
  wire [0:0] s_6;
  wire [31:0] s_7;
  wire [30:0] s_8;
  wire [31:0] s_9;
  wire [31:0] s_10;
  wire [31:0] s_11;
  wire [30:0] s_12;
  wire [31:0] s_13;
  wire [31:0] s_14;
  wire [31:0] s_15;
  wire [30:0] s_16;
  wire [31:0] s_17;
  wire [31:0] s_18;
  wire [8:0] s_19;
  wire [8:0] s_20;
  wire [7:0] s_21;
  wire [22:0] s_22;
  wire [23:0] s_23;
  wire [0:0] s_24;
  wire [23:0] s_25;
  wire [23:0] s_26;
  wire [23:0] s_27;
  wire [24:0] s_28;
  wire [24:0] s_29;
  wire [24:0] s_30;
  wire [24:0] s_31;
  wire [23:0] s_32;
  wire [26:0] s_33;
  wire [26:0] s_34;
  wire [26:0] s_35;
  wire [26:0] s_36;
  wire [26:0] s_37;
  wire [26:0] s_38;
  wire [26:0] s_39;
  wire [26:0] s_40;
  wire [26:0] s_41;
  wire [26:0] s_42;
  wire [26:0] s_43;
  wire [26:0] s_44;
  wire [26:0] s_45;
  wire [26:0] s_46;
  wire [26:0] s_47;
  wire [26:0] s_48;
  wire [26:0] s_49;
  wire [26:0] s_50;
  wire [26:0] s_51;
  wire [26:0] s_52;
  wire [26:0] s_53;
  wire [26:0] s_54;
  wire [26:0] s_55;
  wire [26:0] s_56;
  wire [26:0] s_57;
  wire [26:0] s_58;
  wire [26:0] s_59;
  wire [26:0] s_60;
  wire [26:0] s_61;
  wire [26:0] s_62;
  wire [26:0] s_63;
  wire [26:0] s_64;
  wire [26:0] s_65;
  wire [26:0] s_66;
  wire [26:0] s_67;
  wire [26:0] s_68;
  wire [26:0] s_69;
  wire [26:0] s_70;
  wire [26:0] s_71;
  wire [26:0] s_72;
  wire [26:0] s_73;
  wire [26:0] s_74;
  wire [26:0] s_75;
  wire [26:0] s_76;
  wire [26:0] s_77;
  wire [26:0] s_78;
  wire [26:0] s_79;
  wire [26:0] s_80;
  wire [26:0] s_81;
  wire [26:0] s_82;
  wire [26:0] s_83;
  wire [26:0] s_84;
  wire [26:0] s_85;
  wire [26:0] s_86;
  wire [26:0] s_87;
  wire [26:0] s_88;
  wire [26:0] s_89;
  wire [26:0] s_90;
  wire [26:0] s_91;
  wire [26:0] s_92;
  wire [26:0] s_93;
  wire [26:0] s_94;
  wire [26:0] s_95;
  wire [26:0] s_96;
  wire [26:0] s_97;
  wire [26:0] s_98;
  wire [26:0] s_99;
  wire [26:0] s_100;
  wire [26:0] s_101;
  wire [26:0] s_102;
  wire [26:0] s_103;
  wire [26:0] s_104;
  wire [26:0] s_105;
  wire [26:0] s_106;
  wire [26:0] s_107;
  wire [26:0] s_108;
  wire [26:0] s_109;
  wire [26:0] s_110;
  wire [26:0] s_111;
  wire [26:0] s_112;
  wire [26:0] s_113;
  wire [26:0] s_114;
  wire [26:0] s_115;
  wire [26:0] s_116;
  wire [26:0] s_117;
  wire [26:0] s_118;
  wire [26:0] s_119;
  wire [26:0] s_120;
  wire [26:0] s_121;
  wire [0:0] s_122;
  wire [26:0] s_123;
  wire [26:0] s_124;
  wire [0:0] s_125;
  wire [0:0] s_126;
  wire [27:0] s_127;
  wire [27:0] s_128;
  wire [26:0] s_129;
  wire [26:0] s_130;
  wire [23:0] s_131;
  wire [23:0] s_132;
  wire [23:0] s_133;
  wire [23:0] s_134;
  wire [0:0] s_135;
  wire [0:0] s_136;
  wire [0:0] s_137;
  wire [0:0] s_138;
  wire [7:0] s_139;
  wire [7:0] s_140;
  wire [6:0] s_141;
  wire [7:0] s_142;
  wire [22:0] s_143;
  wire [9:0] s_144;
  wire [9:0] s_145;
  wire [5:0] s_146;
  wire [5:0] s_147;
  wire [0:0] s_148;
  wire [0:0] s_149;
  wire [4:0] s_150;
  wire [0:0] s_151;
  wire [0:0] s_152;
  wire [3:0] s_153;
  wire [0:0] s_154;
  wire [0:0] s_155;
  wire [2:0] s_156;
  wire [0:0] s_157;
  wire [0:0] s_158;
  wire [1:0] s_159;
  wire [0:0] s_160;
  wire [0:0] s_161;
  wire [0:0] s_162;
  wire [1:0] s_163;
  wire [3:0] s_164;
  wire [7:0] s_165;
  wire [15:0] s_166;
  wire [31:0] s_167;
  wire [30:0] s_168;
  wire [29:0] s_169;
  wire [28:0] s_170;
  wire [27:0] s_171;
  wire [26:0] s_172;
  wire [25:0] s_173;
  wire [24:0] s_174;
  wire [0:0] s_175;
  wire [0:0] s_176;
  wire [0:0] s_177;
  wire [0:0] s_178;
  wire [0:0] s_179;
  wire [0:0] s_180;
  wire [0:0] s_181;
  wire [0:0] s_182;
  wire [0:0] s_183;
  wire [0:0] s_184;
  wire [0:0] s_185;
  wire [0:0] s_186;
  wire [0:0] s_187;
  wire [0:0] s_188;
  wire [0:0] s_189;
  wire [1:0] s_190;
  wire [0:0] s_191;
  wire [0:0] s_192;
  wire [0:0] s_193;
  wire [1:0] s_194;
  wire [0:0] s_195;
  wire [0:0] s_196;
  wire [0:0] s_197;
  wire [0:0] s_198;
  wire [0:0] s_199;
  wire [0:0] s_200;
  wire [1:0] s_201;
  wire [0:0] s_202;
  wire [0:0] s_203;
  wire [0:0] s_204;
  wire [0:0] s_205;
  wire [0:0] s_206;
  wire [0:0] s_207;
  wire [2:0] s_208;
  wire [0:0] s_209;
  wire [0:0] s_210;
  wire [1:0] s_211;
  wire [0:0] s_212;
  wire [0:0] s_213;
  wire [0:0] s_214;
  wire [1:0] s_215;
  wire [3:0] s_216;
  wire [0:0] s_217;
  wire [0:0] s_218;
  wire [0:0] s_219;
  wire [0:0] s_220;
  wire [0:0] s_221;
  wire [0:0] s_222;
  wire [0:0] s_223;
  wire [1:0] s_224;
  wire [0:0] s_225;
  wire [0:0] s_226;
  wire [0:0] s_227;
  wire [1:0] s_228;
  wire [0:0] s_229;
  wire [0:0] s_230;
  wire [0:0] s_231;
  wire [0:0] s_232;
  wire [0:0] s_233;
  wire [0:0] s_234;
  wire [1:0] s_235;
  wire [0:0] s_236;
  wire [0:0] s_237;
  wire [0:0] s_238;
  wire [0:0] s_239;
  wire [0:0] s_240;
  wire [2:0] s_241;
  wire [0:0] s_242;
  wire [0:0] s_243;
  wire [1:0] s_244;
  wire [1:0] s_245;
  wire [1:0] s_246;
  wire [0:0] s_247;
  wire [3:0] s_248;
  wire [0:0] s_249;
  wire [0:0] s_250;
  wire [2:0] s_251;
  wire [0:0] s_252;
  wire [0:0] s_253;
  wire [1:0] s_254;
  wire [0:0] s_255;
  wire [0:0] s_256;
  wire [0:0] s_257;
  wire [1:0] s_258;
  wire [3:0] s_259;
  wire [7:0] s_260;
  wire [0:0] s_261;
  wire [0:0] s_262;
  wire [0:0] s_263;
  wire [0:0] s_264;
  wire [0:0] s_265;
  wire [0:0] s_266;
  wire [0:0] s_267;
  wire [1:0] s_268;
  wire [0:0] s_269;
  wire [0:0] s_270;
  wire [0:0] s_271;
  wire [1:0] s_272;
  wire [0:0] s_273;
  wire [0:0] s_274;
  wire [0:0] s_275;
  wire [0:0] s_276;
  wire [0:0] s_277;
  wire [0:0] s_278;
  wire [1:0] s_279;
  wire [0:0] s_280;
  wire [0:0] s_281;
  wire [0:0] s_282;
  wire [0:0] s_283;
  wire [0:0] s_284;
  wire [0:0] s_285;
  wire [2:0] s_286;
  wire [0:0] s_287;
  wire [0:0] s_288;
  wire [1:0] s_289;
  wire [0:0] s_290;
  wire [0:0] s_291;
  wire [0:0] s_292;
  wire [1:0] s_293;
  wire [3:0] s_294;
  wire [0:0] s_295;
  wire [0:0] s_296;
  wire [0:0] s_297;
  wire [0:0] s_298;
  wire [0:0] s_299;
  wire [0:0] s_300;
  wire [0:0] s_301;
  wire [1:0] s_302;
  wire [0:0] s_303;
  wire [0:0] s_304;
  wire [0:0] s_305;
  wire [1:0] s_306;
  wire [0:0] s_307;
  wire [0:0] s_308;
  wire [0:0] s_309;
  wire [0:0] s_310;
  wire [0:0] s_311;
  wire [0:0] s_312;
  wire [1:0] s_313;
  wire [0:0] s_314;
  wire [0:0] s_315;
  wire [0:0] s_316;
  wire [0:0] s_317;
  wire [0:0] s_318;
  wire [2:0] s_319;
  wire [0:0] s_320;
  wire [0:0] s_321;
  wire [1:0] s_322;
  wire [1:0] s_323;
  wire [1:0] s_324;
  wire [3:0] s_325;
  wire [0:0] s_326;
  wire [0:0] s_327;
  wire [2:0] s_328;
  wire [2:0] s_329;
  wire [2:0] s_330;
  wire [0:0] s_331;
  wire [4:0] s_332;
  wire [0:0] s_333;
  wire [0:0] s_334;
  wire [3:0] s_335;
  wire [0:0] s_336;
  wire [0:0] s_337;
  wire [2:0] s_338;
  wire [0:0] s_339;
  wire [0:0] s_340;
  wire [1:0] s_341;
  wire [0:0] s_342;
  wire [0:0] s_343;
  wire [0:0] s_344;
  wire [1:0] s_345;
  wire [3:0] s_346;
  wire [7:0] s_347;
  wire [15:0] s_348;
  wire [0:0] s_349;
  wire [0:0] s_350;
  wire [0:0] s_351;
  wire [0:0] s_352;
  wire [0:0] s_353;
  wire [0:0] s_354;
  wire [0:0] s_355;
  wire [1:0] s_356;
  wire [0:0] s_357;
  wire [0:0] s_358;
  wire [0:0] s_359;
  wire [1:0] s_360;
  wire [0:0] s_361;
  wire [0:0] s_362;
  wire [0:0] s_363;
  wire [0:0] s_364;
  wire [0:0] s_365;
  wire [0:0] s_366;
  wire [1:0] s_367;
  wire [0:0] s_368;
  wire [0:0] s_369;
  wire [0:0] s_370;
  wire [0:0] s_371;
  wire [0:0] s_372;
  wire [0:0] s_373;
  wire [2:0] s_374;
  wire [0:0] s_375;
  wire [0:0] s_376;
  wire [1:0] s_377;
  wire [0:0] s_378;
  wire [0:0] s_379;
  wire [0:0] s_380;
  wire [1:0] s_381;
  wire [3:0] s_382;
  wire [0:0] s_383;
  wire [0:0] s_384;
  wire [0:0] s_385;
  wire [0:0] s_386;
  wire [0:0] s_387;
  wire [0:0] s_388;
  wire [0:0] s_389;
  wire [1:0] s_390;
  wire [0:0] s_391;
  wire [0:0] s_392;
  wire [0:0] s_393;
  wire [1:0] s_394;
  wire [0:0] s_395;
  wire [0:0] s_396;
  wire [0:0] s_397;
  wire [0:0] s_398;
  wire [0:0] s_399;
  wire [0:0] s_400;
  wire [1:0] s_401;
  wire [0:0] s_402;
  wire [0:0] s_403;
  wire [0:0] s_404;
  wire [0:0] s_405;
  wire [0:0] s_406;
  wire [2:0] s_407;
  wire [0:0] s_408;
  wire [0:0] s_409;
  wire [1:0] s_410;
  wire [1:0] s_411;
  wire [1:0] s_412;
  wire [0:0] s_413;
  wire [3:0] s_414;
  wire [0:0] s_415;
  wire [0:0] s_416;
  wire [2:0] s_417;
  wire [0:0] s_418;
  wire [0:0] s_419;
  wire [1:0] s_420;
  wire [0:0] s_421;
  wire [0:0] s_422;
  wire [0:0] s_423;
  wire [1:0] s_424;
  wire [3:0] s_425;
  wire [7:0] s_426;
  wire [0:0] s_427;
  wire [0:0] s_428;
  wire [0:0] s_429;
  wire [0:0] s_430;
  wire [0:0] s_431;
  wire [0:0] s_432;
  wire [0:0] s_433;
  wire [1:0] s_434;
  wire [0:0] s_435;
  wire [0:0] s_436;
  wire [0:0] s_437;
  wire [1:0] s_438;
  wire [0:0] s_439;
  wire [0:0] s_440;
  wire [0:0] s_441;
  wire [0:0] s_442;
  wire [0:0] s_443;
  wire [0:0] s_444;
  wire [1:0] s_445;
  wire [0:0] s_446;
  wire [0:0] s_447;
  wire [0:0] s_448;
  wire [0:0] s_449;
  wire [0:0] s_450;
  wire [0:0] s_451;
  wire [2:0] s_452;
  wire [0:0] s_453;
  wire [0:0] s_454;
  wire [1:0] s_455;
  wire [0:0] s_456;
  wire [0:0] s_457;
  wire [0:0] s_458;
  wire [1:0] s_459;
  wire [3:0] s_460;
  wire [0:0] s_461;
  wire [0:0] s_462;
  wire [0:0] s_463;
  wire [0:0] s_464;
  wire [0:0] s_465;
  wire [0:0] s_466;
  wire [0:0] s_467;
  wire [1:0] s_468;
  wire [0:0] s_469;
  wire [0:0] s_470;
  wire [0:0] s_471;
  wire [1:0] s_472;
  wire [0:0] s_473;
  wire [0:0] s_474;
  wire [0:0] s_475;
  wire [0:0] s_476;
  wire [0:0] s_477;
  wire [0:0] s_478;
  wire [1:0] s_479;
  wire [0:0] s_480;
  wire [0:0] s_481;
  wire [0:0] s_482;
  wire [0:0] s_483;
  wire [0:0] s_484;
  wire [2:0] s_485;
  wire [0:0] s_486;
  wire [0:0] s_487;
  wire [1:0] s_488;
  wire [1:0] s_489;
  wire [1:0] s_490;
  wire [3:0] s_491;
  wire [0:0] s_492;
  wire [0:0] s_493;
  wire [2:0] s_494;
  wire [2:0] s_495;
  wire [2:0] s_496;
  wire [4:0] s_497;
  wire [0:0] s_498;
  wire [0:0] s_499;
  wire [3:0] s_500;
  wire [3:0] s_501;
  wire [3:0] s_502;
  wire [9:0] s_503;
  wire [9:0] s_504;
  wire [9:0] s_505;
  wire [7:0] s_506;
  wire [7:0] s_507;
  wire [9:0] s_508;
  wire [0:0] s_509;
  wire [9:0] s_510;
  wire [9:0] s_511;
  wire [1:0] s_512;
  wire [26:0] s_513;
  wire [26:0] s_514;
  wire [23:0] s_515;
  wire [23:0] s_516;
  wire [23:0] s_517;
  wire [23:0] s_518;
  wire [0:0] s_519;
  wire [0:0] s_520;
  wire [0:0] s_521;
  wire [0:0] s_522;
  wire [7:0] s_523;
  wire [7:0] s_524;
  wire [6:0] s_525;
  wire [7:0] s_526;
  wire [22:0] s_527;
  wire [9:0] s_528;
  wire [9:0] s_529;
  wire [5:0] s_530;
  wire [5:0] s_531;
  wire [0:0] s_532;
  wire [0:0] s_533;
  wire [4:0] s_534;
  wire [0:0] s_535;
  wire [0:0] s_536;
  wire [3:0] s_537;
  wire [0:0] s_538;
  wire [0:0] s_539;
  wire [2:0] s_540;
  wire [0:0] s_541;
  wire [0:0] s_542;
  wire [1:0] s_543;
  wire [0:0] s_544;
  wire [0:0] s_545;
  wire [0:0] s_546;
  wire [1:0] s_547;
  wire [3:0] s_548;
  wire [7:0] s_549;
  wire [15:0] s_550;
  wire [31:0] s_551;
  wire [30:0] s_552;
  wire [29:0] s_553;
  wire [28:0] s_554;
  wire [27:0] s_555;
  wire [26:0] s_556;
  wire [25:0] s_557;
  wire [24:0] s_558;
  wire [0:0] s_559;
  wire [0:0] s_560;
  wire [0:0] s_561;
  wire [0:0] s_562;
  wire [0:0] s_563;
  wire [0:0] s_564;
  wire [0:0] s_565;
  wire [0:0] s_566;
  wire [0:0] s_567;
  wire [0:0] s_568;
  wire [0:0] s_569;
  wire [0:0] s_570;
  wire [0:0] s_571;
  wire [0:0] s_572;
  wire [0:0] s_573;
  wire [1:0] s_574;
  wire [0:0] s_575;
  wire [0:0] s_576;
  wire [0:0] s_577;
  wire [1:0] s_578;
  wire [0:0] s_579;
  wire [0:0] s_580;
  wire [0:0] s_581;
  wire [0:0] s_582;
  wire [0:0] s_583;
  wire [0:0] s_584;
  wire [1:0] s_585;
  wire [0:0] s_586;
  wire [0:0] s_587;
  wire [0:0] s_588;
  wire [0:0] s_589;
  wire [0:0] s_590;
  wire [0:0] s_591;
  wire [2:0] s_592;
  wire [0:0] s_593;
  wire [0:0] s_594;
  wire [1:0] s_595;
  wire [0:0] s_596;
  wire [0:0] s_597;
  wire [0:0] s_598;
  wire [1:0] s_599;
  wire [3:0] s_600;
  wire [0:0] s_601;
  wire [0:0] s_602;
  wire [0:0] s_603;
  wire [0:0] s_604;
  wire [0:0] s_605;
  wire [0:0] s_606;
  wire [0:0] s_607;
  wire [1:0] s_608;
  wire [0:0] s_609;
  wire [0:0] s_610;
  wire [0:0] s_611;
  wire [1:0] s_612;
  wire [0:0] s_613;
  wire [0:0] s_614;
  wire [0:0] s_615;
  wire [0:0] s_616;
  wire [0:0] s_617;
  wire [0:0] s_618;
  wire [1:0] s_619;
  wire [0:0] s_620;
  wire [0:0] s_621;
  wire [0:0] s_622;
  wire [0:0] s_623;
  wire [0:0] s_624;
  wire [2:0] s_625;
  wire [0:0] s_626;
  wire [0:0] s_627;
  wire [1:0] s_628;
  wire [1:0] s_629;
  wire [1:0] s_630;
  wire [0:0] s_631;
  wire [3:0] s_632;
  wire [0:0] s_633;
  wire [0:0] s_634;
  wire [2:0] s_635;
  wire [0:0] s_636;
  wire [0:0] s_637;
  wire [1:0] s_638;
  wire [0:0] s_639;
  wire [0:0] s_640;
  wire [0:0] s_641;
  wire [1:0] s_642;
  wire [3:0] s_643;
  wire [7:0] s_644;
  wire [0:0] s_645;
  wire [0:0] s_646;
  wire [0:0] s_647;
  wire [0:0] s_648;
  wire [0:0] s_649;
  wire [0:0] s_650;
  wire [0:0] s_651;
  wire [1:0] s_652;
  wire [0:0] s_653;
  wire [0:0] s_654;
  wire [0:0] s_655;
  wire [1:0] s_656;
  wire [0:0] s_657;
  wire [0:0] s_658;
  wire [0:0] s_659;
  wire [0:0] s_660;
  wire [0:0] s_661;
  wire [0:0] s_662;
  wire [1:0] s_663;
  wire [0:0] s_664;
  wire [0:0] s_665;
  wire [0:0] s_666;
  wire [0:0] s_667;
  wire [0:0] s_668;
  wire [0:0] s_669;
  wire [2:0] s_670;
  wire [0:0] s_671;
  wire [0:0] s_672;
  wire [1:0] s_673;
  wire [0:0] s_674;
  wire [0:0] s_675;
  wire [0:0] s_676;
  wire [1:0] s_677;
  wire [3:0] s_678;
  wire [0:0] s_679;
  wire [0:0] s_680;
  wire [0:0] s_681;
  wire [0:0] s_682;
  wire [0:0] s_683;
  wire [0:0] s_684;
  wire [0:0] s_685;
  wire [1:0] s_686;
  wire [0:0] s_687;
  wire [0:0] s_688;
  wire [0:0] s_689;
  wire [1:0] s_690;
  wire [0:0] s_691;
  wire [0:0] s_692;
  wire [0:0] s_693;
  wire [0:0] s_694;
  wire [0:0] s_695;
  wire [0:0] s_696;
  wire [1:0] s_697;
  wire [0:0] s_698;
  wire [0:0] s_699;
  wire [0:0] s_700;
  wire [0:0] s_701;
  wire [0:0] s_702;
  wire [2:0] s_703;
  wire [0:0] s_704;
  wire [0:0] s_705;
  wire [1:0] s_706;
  wire [1:0] s_707;
  wire [1:0] s_708;
  wire [3:0] s_709;
  wire [0:0] s_710;
  wire [0:0] s_711;
  wire [2:0] s_712;
  wire [2:0] s_713;
  wire [2:0] s_714;
  wire [0:0] s_715;
  wire [4:0] s_716;
  wire [0:0] s_717;
  wire [0:0] s_718;
  wire [3:0] s_719;
  wire [0:0] s_720;
  wire [0:0] s_721;
  wire [2:0] s_722;
  wire [0:0] s_723;
  wire [0:0] s_724;
  wire [1:0] s_725;
  wire [0:0] s_726;
  wire [0:0] s_727;
  wire [0:0] s_728;
  wire [1:0] s_729;
  wire [3:0] s_730;
  wire [7:0] s_731;
  wire [15:0] s_732;
  wire [0:0] s_733;
  wire [0:0] s_734;
  wire [0:0] s_735;
  wire [0:0] s_736;
  wire [0:0] s_737;
  wire [0:0] s_738;
  wire [0:0] s_739;
  wire [1:0] s_740;
  wire [0:0] s_741;
  wire [0:0] s_742;
  wire [0:0] s_743;
  wire [1:0] s_744;
  wire [0:0] s_745;
  wire [0:0] s_746;
  wire [0:0] s_747;
  wire [0:0] s_748;
  wire [0:0] s_749;
  wire [0:0] s_750;
  wire [1:0] s_751;
  wire [0:0] s_752;
  wire [0:0] s_753;
  wire [0:0] s_754;
  wire [0:0] s_755;
  wire [0:0] s_756;
  wire [0:0] s_757;
  wire [2:0] s_758;
  wire [0:0] s_759;
  wire [0:0] s_760;
  wire [1:0] s_761;
  wire [0:0] s_762;
  wire [0:0] s_763;
  wire [0:0] s_764;
  wire [1:0] s_765;
  wire [3:0] s_766;
  wire [0:0] s_767;
  wire [0:0] s_768;
  wire [0:0] s_769;
  wire [0:0] s_770;
  wire [0:0] s_771;
  wire [0:0] s_772;
  wire [0:0] s_773;
  wire [1:0] s_774;
  wire [0:0] s_775;
  wire [0:0] s_776;
  wire [0:0] s_777;
  wire [1:0] s_778;
  wire [0:0] s_779;
  wire [0:0] s_780;
  wire [0:0] s_781;
  wire [0:0] s_782;
  wire [0:0] s_783;
  wire [0:0] s_784;
  wire [1:0] s_785;
  wire [0:0] s_786;
  wire [0:0] s_787;
  wire [0:0] s_788;
  wire [0:0] s_789;
  wire [0:0] s_790;
  wire [2:0] s_791;
  wire [0:0] s_792;
  wire [0:0] s_793;
  wire [1:0] s_794;
  wire [1:0] s_795;
  wire [1:0] s_796;
  wire [0:0] s_797;
  wire [3:0] s_798;
  wire [0:0] s_799;
  wire [0:0] s_800;
  wire [2:0] s_801;
  wire [0:0] s_802;
  wire [0:0] s_803;
  wire [1:0] s_804;
  wire [0:0] s_805;
  wire [0:0] s_806;
  wire [0:0] s_807;
  wire [1:0] s_808;
  wire [3:0] s_809;
  wire [7:0] s_810;
  wire [0:0] s_811;
  wire [0:0] s_812;
  wire [0:0] s_813;
  wire [0:0] s_814;
  wire [0:0] s_815;
  wire [0:0] s_816;
  wire [0:0] s_817;
  wire [1:0] s_818;
  wire [0:0] s_819;
  wire [0:0] s_820;
  wire [0:0] s_821;
  wire [1:0] s_822;
  wire [0:0] s_823;
  wire [0:0] s_824;
  wire [0:0] s_825;
  wire [0:0] s_826;
  wire [0:0] s_827;
  wire [0:0] s_828;
  wire [1:0] s_829;
  wire [0:0] s_830;
  wire [0:0] s_831;
  wire [0:0] s_832;
  wire [0:0] s_833;
  wire [0:0] s_834;
  wire [0:0] s_835;
  wire [2:0] s_836;
  wire [0:0] s_837;
  wire [0:0] s_838;
  wire [1:0] s_839;
  wire [0:0] s_840;
  wire [0:0] s_841;
  wire [0:0] s_842;
  wire [1:0] s_843;
  wire [3:0] s_844;
  wire [0:0] s_845;
  wire [0:0] s_846;
  wire [0:0] s_847;
  wire [0:0] s_848;
  wire [0:0] s_849;
  wire [0:0] s_850;
  wire [0:0] s_851;
  wire [1:0] s_852;
  wire [0:0] s_853;
  wire [0:0] s_854;
  wire [0:0] s_855;
  wire [1:0] s_856;
  wire [0:0] s_857;
  wire [0:0] s_858;
  wire [0:0] s_859;
  wire [0:0] s_860;
  wire [0:0] s_861;
  wire [0:0] s_862;
  wire [1:0] s_863;
  wire [0:0] s_864;
  wire [0:0] s_865;
  wire [0:0] s_866;
  wire [0:0] s_867;
  wire [0:0] s_868;
  wire [2:0] s_869;
  wire [0:0] s_870;
  wire [0:0] s_871;
  wire [1:0] s_872;
  wire [1:0] s_873;
  wire [1:0] s_874;
  wire [3:0] s_875;
  wire [0:0] s_876;
  wire [0:0] s_877;
  wire [2:0] s_878;
  wire [2:0] s_879;
  wire [2:0] s_880;
  wire [4:0] s_881;
  wire [0:0] s_882;
  wire [0:0] s_883;
  wire [3:0] s_884;
  wire [3:0] s_885;
  wire [3:0] s_886;
  wire [9:0] s_887;
  wire [9:0] s_888;
  wire [9:0] s_889;
  wire [7:0] s_890;
  wire [7:0] s_891;
  wire [9:0] s_892;
  wire [0:0] s_893;
  wire [9:0] s_894;
  wire [9:0] s_895;
  wire [1:0] s_896;
  wire [0:0] s_897;
  wire [26:0] s_898;
  wire [0:0] s_899;
  wire [0:0] s_900;
  wire [27:0] s_901;
  wire [27:0] s_902;
  wire [27:0] s_903;
  wire [27:0] s_904;
  wire [27:0] s_905;
  wire [27:0] s_906;
  wire [0:0] s_907;
  wire [0:0] s_908;
  wire [26:0] s_909;
  wire [0:0] s_910;
  wire [26:0] s_911;
  wire [0:0] s_912;
  wire [0:0] s_913;
  wire [27:0] s_914;
  wire [27:0] s_915;
  wire [27:0] s_916;
  wire [27:0] s_917;
  wire [27:0] s_918;
  wire [27:0] s_919;
  wire [0:0] s_920;
  wire [0:0] s_921;
  wire [26:0] s_922;
  wire [0:0] s_923;
  wire [26:0] s_924;
  wire [0:0] s_925;
  wire [0:0] s_926;
  wire [27:0] s_927;
  wire [27:0] s_928;
  wire [27:0] s_929;
  wire [27:0] s_930;
  wire [27:0] s_931;
  wire [27:0] s_932;
  wire [0:0] s_933;
  wire [0:0] s_934;
  wire [26:0] s_935;
  wire [0:0] s_936;
  wire [26:0] s_937;
  wire [0:0] s_938;
  wire [0:0] s_939;
  wire [27:0] s_940;
  wire [27:0] s_941;
  wire [27:0] s_942;
  wire [27:0] s_943;
  wire [27:0] s_944;
  wire [27:0] s_945;
  wire [0:0] s_946;
  wire [0:0] s_947;
  wire [26:0] s_948;
  wire [0:0] s_949;
  wire [26:0] s_950;
  wire [0:0] s_951;
  wire [0:0] s_952;
  wire [27:0] s_953;
  wire [27:0] s_954;
  wire [27:0] s_955;
  wire [27:0] s_956;
  wire [27:0] s_957;
  wire [27:0] s_958;
  wire [0:0] s_959;
  wire [0:0] s_960;
  wire [26:0] s_961;
  wire [0:0] s_962;
  wire [26:0] s_963;
  wire [0:0] s_964;
  wire [0:0] s_965;
  wire [27:0] s_966;
  wire [27:0] s_967;
  wire [27:0] s_968;
  wire [27:0] s_969;
  wire [27:0] s_970;
  wire [27:0] s_971;
  wire [0:0] s_972;
  wire [0:0] s_973;
  wire [26:0] s_974;
  wire [0:0] s_975;
  wire [26:0] s_976;
  wire [0:0] s_977;
  wire [0:0] s_978;
  wire [27:0] s_979;
  wire [27:0] s_980;
  wire [27:0] s_981;
  wire [27:0] s_982;
  wire [27:0] s_983;
  wire [27:0] s_984;
  wire [0:0] s_985;
  wire [0:0] s_986;
  wire [26:0] s_987;
  wire [0:0] s_988;
  wire [26:0] s_989;
  wire [0:0] s_990;
  wire [0:0] s_991;
  wire [27:0] s_992;
  wire [27:0] s_993;
  wire [27:0] s_994;
  wire [27:0] s_995;
  wire [27:0] s_996;
  wire [27:0] s_997;
  wire [0:0] s_998;
  wire [0:0] s_999;
  wire [26:0] s_1000;
  wire [0:0] s_1001;
  wire [26:0] s_1002;
  wire [0:0] s_1003;
  wire [0:0] s_1004;
  wire [27:0] s_1005;
  wire [27:0] s_1006;
  wire [27:0] s_1007;
  wire [27:0] s_1008;
  wire [27:0] s_1009;
  wire [27:0] s_1010;
  wire [0:0] s_1011;
  wire [0:0] s_1012;
  wire [26:0] s_1013;
  wire [0:0] s_1014;
  wire [26:0] s_1015;
  wire [0:0] s_1016;
  wire [0:0] s_1017;
  wire [27:0] s_1018;
  wire [27:0] s_1019;
  wire [27:0] s_1020;
  wire [27:0] s_1021;
  wire [27:0] s_1022;
  wire [27:0] s_1023;
  wire [0:0] s_1024;
  wire [0:0] s_1025;
  wire [26:0] s_1026;
  wire [0:0] s_1027;
  wire [26:0] s_1028;
  wire [0:0] s_1029;
  wire [0:0] s_1030;
  wire [27:0] s_1031;
  wire [27:0] s_1032;
  wire [27:0] s_1033;
  wire [27:0] s_1034;
  wire [27:0] s_1035;
  wire [27:0] s_1036;
  wire [0:0] s_1037;
  wire [0:0] s_1038;
  wire [26:0] s_1039;
  wire [0:0] s_1040;
  wire [26:0] s_1041;
  wire [0:0] s_1042;
  wire [0:0] s_1043;
  wire [27:0] s_1044;
  wire [27:0] s_1045;
  wire [27:0] s_1046;
  wire [27:0] s_1047;
  wire [27:0] s_1048;
  wire [27:0] s_1049;
  wire [0:0] s_1050;
  wire [0:0] s_1051;
  wire [26:0] s_1052;
  wire [0:0] s_1053;
  wire [26:0] s_1054;
  wire [0:0] s_1055;
  wire [0:0] s_1056;
  wire [27:0] s_1057;
  wire [27:0] s_1058;
  wire [27:0] s_1059;
  wire [27:0] s_1060;
  wire [27:0] s_1061;
  wire [27:0] s_1062;
  wire [0:0] s_1063;
  wire [0:0] s_1064;
  wire [26:0] s_1065;
  wire [0:0] s_1066;
  wire [26:0] s_1067;
  wire [0:0] s_1068;
  wire [0:0] s_1069;
  wire [27:0] s_1070;
  wire [27:0] s_1071;
  wire [27:0] s_1072;
  wire [27:0] s_1073;
  wire [27:0] s_1074;
  wire [27:0] s_1075;
  wire [0:0] s_1076;
  wire [0:0] s_1077;
  wire [26:0] s_1078;
  wire [0:0] s_1079;
  wire [26:0] s_1080;
  wire [0:0] s_1081;
  wire [0:0] s_1082;
  wire [27:0] s_1083;
  wire [27:0] s_1084;
  wire [27:0] s_1085;
  wire [27:0] s_1086;
  wire [27:0] s_1087;
  wire [27:0] s_1088;
  wire [0:0] s_1089;
  wire [0:0] s_1090;
  wire [26:0] s_1091;
  wire [0:0] s_1092;
  wire [26:0] s_1093;
  wire [0:0] s_1094;
  wire [0:0] s_1095;
  wire [27:0] s_1096;
  wire [27:0] s_1097;
  wire [27:0] s_1098;
  wire [27:0] s_1099;
  wire [27:0] s_1100;
  wire [27:0] s_1101;
  wire [0:0] s_1102;
  wire [0:0] s_1103;
  wire [26:0] s_1104;
  wire [0:0] s_1105;
  wire [26:0] s_1106;
  wire [0:0] s_1107;
  wire [0:0] s_1108;
  wire [27:0] s_1109;
  wire [27:0] s_1110;
  wire [27:0] s_1111;
  wire [27:0] s_1112;
  wire [27:0] s_1113;
  wire [27:0] s_1114;
  wire [0:0] s_1115;
  wire [0:0] s_1116;
  wire [26:0] s_1117;
  wire [0:0] s_1118;
  wire [26:0] s_1119;
  wire [0:0] s_1120;
  wire [0:0] s_1121;
  wire [27:0] s_1122;
  wire [27:0] s_1123;
  wire [27:0] s_1124;
  wire [27:0] s_1125;
  wire [27:0] s_1126;
  wire [27:0] s_1127;
  wire [0:0] s_1128;
  wire [0:0] s_1129;
  wire [26:0] s_1130;
  wire [0:0] s_1131;
  wire [26:0] s_1132;
  wire [0:0] s_1133;
  wire [0:0] s_1134;
  wire [27:0] s_1135;
  wire [27:0] s_1136;
  wire [27:0] s_1137;
  wire [27:0] s_1138;
  wire [27:0] s_1139;
  wire [27:0] s_1140;
  wire [0:0] s_1141;
  wire [0:0] s_1142;
  wire [26:0] s_1143;
  wire [0:0] s_1144;
  wire [26:0] s_1145;
  wire [0:0] s_1146;
  wire [0:0] s_1147;
  wire [27:0] s_1148;
  wire [27:0] s_1149;
  wire [27:0] s_1150;
  wire [27:0] s_1151;
  wire [27:0] s_1152;
  wire [27:0] s_1153;
  wire [0:0] s_1154;
  wire [0:0] s_1155;
  wire [26:0] s_1156;
  wire [0:0] s_1157;
  wire [26:0] s_1158;
  wire [0:0] s_1159;
  wire [0:0] s_1160;
  wire [27:0] s_1161;
  wire [27:0] s_1162;
  wire [27:0] s_1163;
  wire [27:0] s_1164;
  wire [27:0] s_1165;
  wire [27:0] s_1166;
  wire [0:0] s_1167;
  wire [0:0] s_1168;
  wire [26:0] s_1169;
  wire [0:0] s_1170;
  wire [26:0] s_1171;
  wire [0:0] s_1172;
  wire [0:0] s_1173;
  wire [27:0] s_1174;
  wire [27:0] s_1175;
  wire [27:0] s_1176;
  wire [27:0] s_1177;
  wire [27:0] s_1178;
  wire [27:0] s_1179;
  wire [0:0] s_1180;
  wire [0:0] s_1181;
  wire [26:0] s_1182;
  wire [0:0] s_1183;
  wire [26:0] s_1184;
  wire [0:0] s_1185;
  wire [0:0] s_1186;
  wire [27:0] s_1187;
  wire [27:0] s_1188;
  wire [27:0] s_1189;
  wire [27:0] s_1190;
  wire [27:0] s_1191;
  wire [27:0] s_1192;
  wire [0:0] s_1193;
  wire [0:0] s_1194;
  wire [26:0] s_1195;
  wire [0:0] s_1196;
  wire [26:0] s_1197;
  wire [0:0] s_1198;
  wire [0:0] s_1199;
  wire [27:0] s_1200;
  wire [27:0] s_1201;
  wire [27:0] s_1202;
  wire [27:0] s_1203;
  wire [27:0] s_1204;
  wire [27:0] s_1205;
  wire [0:0] s_1206;
  wire [0:0] s_1207;
  wire [26:0] s_1208;
  wire [0:0] s_1209;
  wire [26:0] s_1210;
  wire [0:0] s_1211;
  wire [0:0] s_1212;
  wire [27:0] s_1213;
  wire [27:0] s_1214;
  wire [27:0] s_1215;
  wire [27:0] s_1216;
  wire [27:0] s_1217;
  wire [27:0] s_1218;
  wire [0:0] s_1219;
  wire [0:0] s_1220;
  wire [26:0] s_1221;
  wire [0:0] s_1222;
  wire [26:0] s_1223;
  wire [0:0] s_1224;
  wire [0:0] s_1225;
  wire [27:0] s_1226;
  wire [27:0] s_1227;
  wire [27:0] s_1228;
  wire [27:0] s_1229;
  wire [27:0] s_1230;
  wire [27:0] s_1231;
  wire [0:0] s_1232;
  wire [0:0] s_1233;
  wire [26:0] s_1234;
  wire [9:0] s_1235;
  wire [9:0] s_1236;
  wire [9:0] s_1237;
  wire [0:0] s_1238;
  wire [9:0] s_1239;
  wire [9:0] s_1240;
  wire [9:0] s_1241;
  wire [9:0] s_1242;
  wire [9:0] s_1243;
  wire [9:0] s_1244;
  wire [9:0] s_1245;
  wire [9:0] s_1246;
  wire [9:0] s_1247;
  wire [9:0] s_1248;
  wire [9:0] s_1249;
  wire [0:0] s_1250;
  wire [9:0] s_1251;
  wire [9:0] s_1252;
  wire [5:0] s_1253;
  wire [5:0] s_1254;
  wire [0:0] s_1255;
  wire [0:0] s_1256;
  wire [4:0] s_1257;
  wire [0:0] s_1258;
  wire [0:0] s_1259;
  wire [3:0] s_1260;
  wire [0:0] s_1261;
  wire [0:0] s_1262;
  wire [2:0] s_1263;
  wire [0:0] s_1264;
  wire [0:0] s_1265;
  wire [1:0] s_1266;
  wire [0:0] s_1267;
  wire [0:0] s_1268;
  wire [0:0] s_1269;
  wire [1:0] s_1270;
  wire [3:0] s_1271;
  wire [7:0] s_1272;
  wire [15:0] s_1273;
  wire [31:0] s_1274;
  wire [30:0] s_1275;
  wire [29:0] s_1276;
  wire [28:0] s_1277;
  wire [27:0] s_1278;
  wire [0:0] s_1279;
  wire [0:0] s_1280;
  wire [0:0] s_1281;
  wire [0:0] s_1282;
  wire [0:0] s_1283;
  wire [0:0] s_1284;
  wire [0:0] s_1285;
  wire [0:0] s_1286;
  wire [0:0] s_1287;
  wire [0:0] s_1288;
  wire [0:0] s_1289;
  wire [0:0] s_1290;
  wire [1:0] s_1291;
  wire [0:0] s_1292;
  wire [0:0] s_1293;
  wire [0:0] s_1294;
  wire [1:0] s_1295;
  wire [0:0] s_1296;
  wire [0:0] s_1297;
  wire [0:0] s_1298;
  wire [0:0] s_1299;
  wire [0:0] s_1300;
  wire [0:0] s_1301;
  wire [1:0] s_1302;
  wire [0:0] s_1303;
  wire [0:0] s_1304;
  wire [0:0] s_1305;
  wire [0:0] s_1306;
  wire [0:0] s_1307;
  wire [0:0] s_1308;
  wire [2:0] s_1309;
  wire [0:0] s_1310;
  wire [0:0] s_1311;
  wire [1:0] s_1312;
  wire [0:0] s_1313;
  wire [0:0] s_1314;
  wire [0:0] s_1315;
  wire [1:0] s_1316;
  wire [3:0] s_1317;
  wire [0:0] s_1318;
  wire [0:0] s_1319;
  wire [0:0] s_1320;
  wire [0:0] s_1321;
  wire [0:0] s_1322;
  wire [0:0] s_1323;
  wire [0:0] s_1324;
  wire [1:0] s_1325;
  wire [0:0] s_1326;
  wire [0:0] s_1327;
  wire [0:0] s_1328;
  wire [1:0] s_1329;
  wire [0:0] s_1330;
  wire [0:0] s_1331;
  wire [0:0] s_1332;
  wire [0:0] s_1333;
  wire [0:0] s_1334;
  wire [0:0] s_1335;
  wire [1:0] s_1336;
  wire [0:0] s_1337;
  wire [0:0] s_1338;
  wire [0:0] s_1339;
  wire [0:0] s_1340;
  wire [0:0] s_1341;
  wire [2:0] s_1342;
  wire [0:0] s_1343;
  wire [0:0] s_1344;
  wire [1:0] s_1345;
  wire [1:0] s_1346;
  wire [1:0] s_1347;
  wire [0:0] s_1348;
  wire [3:0] s_1349;
  wire [0:0] s_1350;
  wire [0:0] s_1351;
  wire [2:0] s_1352;
  wire [0:0] s_1353;
  wire [0:0] s_1354;
  wire [1:0] s_1355;
  wire [0:0] s_1356;
  wire [0:0] s_1357;
  wire [0:0] s_1358;
  wire [1:0] s_1359;
  wire [3:0] s_1360;
  wire [7:0] s_1361;
  wire [0:0] s_1362;
  wire [0:0] s_1363;
  wire [0:0] s_1364;
  wire [0:0] s_1365;
  wire [0:0] s_1366;
  wire [0:0] s_1367;
  wire [0:0] s_1368;
  wire [1:0] s_1369;
  wire [0:0] s_1370;
  wire [0:0] s_1371;
  wire [0:0] s_1372;
  wire [1:0] s_1373;
  wire [0:0] s_1374;
  wire [0:0] s_1375;
  wire [0:0] s_1376;
  wire [0:0] s_1377;
  wire [0:0] s_1378;
  wire [0:0] s_1379;
  wire [1:0] s_1380;
  wire [0:0] s_1381;
  wire [0:0] s_1382;
  wire [0:0] s_1383;
  wire [0:0] s_1384;
  wire [0:0] s_1385;
  wire [0:0] s_1386;
  wire [2:0] s_1387;
  wire [0:0] s_1388;
  wire [0:0] s_1389;
  wire [1:0] s_1390;
  wire [0:0] s_1391;
  wire [0:0] s_1392;
  wire [0:0] s_1393;
  wire [1:0] s_1394;
  wire [3:0] s_1395;
  wire [0:0] s_1396;
  wire [0:0] s_1397;
  wire [0:0] s_1398;
  wire [0:0] s_1399;
  wire [0:0] s_1400;
  wire [0:0] s_1401;
  wire [0:0] s_1402;
  wire [1:0] s_1403;
  wire [0:0] s_1404;
  wire [0:0] s_1405;
  wire [0:0] s_1406;
  wire [1:0] s_1407;
  wire [0:0] s_1408;
  wire [0:0] s_1409;
  wire [0:0] s_1410;
  wire [0:0] s_1411;
  wire [0:0] s_1412;
  wire [0:0] s_1413;
  wire [1:0] s_1414;
  wire [0:0] s_1415;
  wire [0:0] s_1416;
  wire [0:0] s_1417;
  wire [0:0] s_1418;
  wire [0:0] s_1419;
  wire [2:0] s_1420;
  wire [0:0] s_1421;
  wire [0:0] s_1422;
  wire [1:0] s_1423;
  wire [1:0] s_1424;
  wire [1:0] s_1425;
  wire [3:0] s_1426;
  wire [0:0] s_1427;
  wire [0:0] s_1428;
  wire [2:0] s_1429;
  wire [2:0] s_1430;
  wire [2:0] s_1431;
  wire [0:0] s_1432;
  wire [4:0] s_1433;
  wire [0:0] s_1434;
  wire [0:0] s_1435;
  wire [3:0] s_1436;
  wire [0:0] s_1437;
  wire [0:0] s_1438;
  wire [2:0] s_1439;
  wire [0:0] s_1440;
  wire [0:0] s_1441;
  wire [1:0] s_1442;
  wire [0:0] s_1443;
  wire [0:0] s_1444;
  wire [0:0] s_1445;
  wire [1:0] s_1446;
  wire [3:0] s_1447;
  wire [7:0] s_1448;
  wire [15:0] s_1449;
  wire [0:0] s_1450;
  wire [0:0] s_1451;
  wire [0:0] s_1452;
  wire [0:0] s_1453;
  wire [0:0] s_1454;
  wire [0:0] s_1455;
  wire [0:0] s_1456;
  wire [1:0] s_1457;
  wire [0:0] s_1458;
  wire [0:0] s_1459;
  wire [0:0] s_1460;
  wire [1:0] s_1461;
  wire [0:0] s_1462;
  wire [0:0] s_1463;
  wire [0:0] s_1464;
  wire [0:0] s_1465;
  wire [0:0] s_1466;
  wire [0:0] s_1467;
  wire [1:0] s_1468;
  wire [0:0] s_1469;
  wire [0:0] s_1470;
  wire [0:0] s_1471;
  wire [0:0] s_1472;
  wire [0:0] s_1473;
  wire [0:0] s_1474;
  wire [2:0] s_1475;
  wire [0:0] s_1476;
  wire [0:0] s_1477;
  wire [1:0] s_1478;
  wire [0:0] s_1479;
  wire [0:0] s_1480;
  wire [0:0] s_1481;
  wire [1:0] s_1482;
  wire [3:0] s_1483;
  wire [0:0] s_1484;
  wire [0:0] s_1485;
  wire [0:0] s_1486;
  wire [0:0] s_1487;
  wire [0:0] s_1488;
  wire [0:0] s_1489;
  wire [0:0] s_1490;
  wire [1:0] s_1491;
  wire [0:0] s_1492;
  wire [0:0] s_1493;
  wire [0:0] s_1494;
  wire [1:0] s_1495;
  wire [0:0] s_1496;
  wire [0:0] s_1497;
  wire [0:0] s_1498;
  wire [0:0] s_1499;
  wire [0:0] s_1500;
  wire [0:0] s_1501;
  wire [1:0] s_1502;
  wire [0:0] s_1503;
  wire [0:0] s_1504;
  wire [0:0] s_1505;
  wire [0:0] s_1506;
  wire [0:0] s_1507;
  wire [2:0] s_1508;
  wire [0:0] s_1509;
  wire [0:0] s_1510;
  wire [1:0] s_1511;
  wire [1:0] s_1512;
  wire [1:0] s_1513;
  wire [0:0] s_1514;
  wire [3:0] s_1515;
  wire [0:0] s_1516;
  wire [0:0] s_1517;
  wire [2:0] s_1518;
  wire [0:0] s_1519;
  wire [0:0] s_1520;
  wire [1:0] s_1521;
  wire [0:0] s_1522;
  wire [0:0] s_1523;
  wire [0:0] s_1524;
  wire [1:0] s_1525;
  wire [3:0] s_1526;
  wire [7:0] s_1527;
  wire [0:0] s_1528;
  wire [0:0] s_1529;
  wire [0:0] s_1530;
  wire [0:0] s_1531;
  wire [0:0] s_1532;
  wire [0:0] s_1533;
  wire [0:0] s_1534;
  wire [1:0] s_1535;
  wire [0:0] s_1536;
  wire [0:0] s_1537;
  wire [0:0] s_1538;
  wire [1:0] s_1539;
  wire [0:0] s_1540;
  wire [0:0] s_1541;
  wire [0:0] s_1542;
  wire [0:0] s_1543;
  wire [0:0] s_1544;
  wire [0:0] s_1545;
  wire [1:0] s_1546;
  wire [0:0] s_1547;
  wire [0:0] s_1548;
  wire [0:0] s_1549;
  wire [0:0] s_1550;
  wire [0:0] s_1551;
  wire [0:0] s_1552;
  wire [2:0] s_1553;
  wire [0:0] s_1554;
  wire [0:0] s_1555;
  wire [1:0] s_1556;
  wire [0:0] s_1557;
  wire [0:0] s_1558;
  wire [0:0] s_1559;
  wire [1:0] s_1560;
  wire [3:0] s_1561;
  wire [0:0] s_1562;
  wire [0:0] s_1563;
  wire [0:0] s_1564;
  wire [0:0] s_1565;
  wire [0:0] s_1566;
  wire [0:0] s_1567;
  wire [0:0] s_1568;
  wire [1:0] s_1569;
  wire [0:0] s_1570;
  wire [0:0] s_1571;
  wire [0:0] s_1572;
  wire [1:0] s_1573;
  wire [0:0] s_1574;
  wire [0:0] s_1575;
  wire [0:0] s_1576;
  wire [0:0] s_1577;
  wire [0:0] s_1578;
  wire [0:0] s_1579;
  wire [1:0] s_1580;
  wire [0:0] s_1581;
  wire [0:0] s_1582;
  wire [0:0] s_1583;
  wire [0:0] s_1584;
  wire [0:0] s_1585;
  wire [2:0] s_1586;
  wire [0:0] s_1587;
  wire [0:0] s_1588;
  wire [1:0] s_1589;
  wire [1:0] s_1590;
  wire [1:0] s_1591;
  wire [3:0] s_1592;
  wire [0:0] s_1593;
  wire [0:0] s_1594;
  wire [2:0] s_1595;
  wire [2:0] s_1596;
  wire [2:0] s_1597;
  wire [4:0] s_1598;
  wire [0:0] s_1599;
  wire [0:0] s_1600;
  wire [3:0] s_1601;
  wire [3:0] s_1602;
  wire [3:0] s_1603;
  wire [9:0] s_1604;
  wire [9:0] s_1605;
  wire [9:0] s_1606;
  wire [9:0] s_1607;
  wire [9:0] s_1608;
  wire [9:0] s_1609;
  wire [0:0] s_1610;
  wire [9:0] s_1611;
  wire [9:0] s_1612;
  wire [1:0] s_1613;
  wire [0:0] s_1614;
  wire [23:0] s_1615;
  wire [0:0] s_1616;
  wire [0:0] s_1617;
  wire [0:0] s_1618;
  wire [0:0] s_1619;
  wire [0:0] s_1620;
  wire [0:0] s_1621;
  wire [0:0] s_1622;
  wire [0:0] s_1623;
  wire [0:0] s_1624;
  wire [0:0] s_1625;
  wire [0:0] s_1626;
  wire [0:0] s_1627;
  wire [27:0] s_1628;
  wire [27:0] s_1629;
  wire [0:0] s_1630;
  wire [0:0] s_1631;
  wire [0:0] s_1632;
  wire [23:0] s_1633;
  wire [0:0] s_1634;
  wire [0:0] s_1635;
  wire [0:0] s_1636;
  wire [0:0] s_1637;
  wire [7:0] s_1638;
  wire [0:0] s_1639;
  wire [22:0] s_1640;
  wire [31:0] s_1641;
  wire [8:0] s_1642;
  wire [0:0] s_1643;
  wire [7:0] s_1644;
  wire [7:0] s_1645;
  wire [9:0] s_1646;
  wire [9:0] s_1647;
  wire [9:0] s_1648;
  wire [9:0] s_1649;
  wire [9:0] s_1650;
  wire [9:0] s_1651;
  wire [6:0] s_1652;
  wire [22:0] s_1653;
  wire [0:0] s_1654;
  wire [0:0] s_1655;
  wire [7:0] s_1656;
  wire [0:0] s_1657;
  wire [0:0] s_1658;
  wire [0:0] s_1659;
  wire [23:0] s_1660;
  wire [0:0] s_1661;
  wire [0:0] s_1662;
  wire [0:0] s_1663;
  wire [0:0] s_1664;
  wire [0:0] s_1665;
  wire [8:0] s_1666;
  wire [0:0] s_1667;
  wire [0:0] s_1668;
  wire [0:0] s_1669;
  wire [7:0] s_1670;
  wire [0:0] s_1671;
  wire [22:0] s_1672;
  wire [0:0] s_1673;
  wire [0:0] s_1674;
  wire [0:0] s_1675;
  wire [0:0] s_1676;
  wire [0:0] s_1677;
  wire [0:0] s_1678;
  wire [0:0] s_1679;
  wire [0:0] s_1680;
  wire [0:0] s_1681;
  wire [0:0] s_1682;
  wire [7:0] s_1683;
  wire [0:0] s_1684;
  wire [22:0] s_1685;
  wire [0:0] s_1686;
  wire [0:0] s_1687;
  wire [7:0] s_1688;
  wire [0:0] s_1689;
  wire [22:0] s_1690;
  wire [0:0] s_1691;

  assign s_0 = s_1678?s_1:s_9;
  dq #(32, 36) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_8};
  assign s_3 = s_4 ^ s_6;
  assign s_4 = s_5[31];
  assign s_5 = div_a;
  assign s_6 = s_7[31];
  assign s_7 = div_b;
  assign s_8 = 31'd2143289344;
  assign s_9 = s_1661?s_10:s_13;
  dq #(32, 36) dq_s_10 (clk, s_10, s_11);
  assign s_11 = {s_3,s_12};
  assign s_12 = 31'd2139095040;
  assign s_13 = s_1659?s_14:s_17;
  dq #(32, 36) dq_s_14 (clk, s_14, s_15);
  assign s_15 = {s_3,s_16};
  assign s_16 = 31'd0;
  assign s_17 = s_1654?s_18:s_1641;
  assign s_18 = {s_19,s_22};
  dq #(9, 36) dq_s_19 (clk, s_19, s_20);
  assign s_20 = {s_3,s_21};
  assign s_21 = 8'd0;
  assign s_22 = s_23[22:0];
  assign s_23 = s_1635?s_24:s_25;
  assign s_24 = 1'd0;
  dq #(24, 1) dq_s_25 (clk, s_25, s_26);
  assign s_26 = s_1634?s_27:s_1633;
  assign s_27 = s_28[24:1];
  assign s_28 = s_1616?s_29:s_1615;
  dq #(25, 1) dq_s_29 (clk, s_29, s_30);
  assign s_30 = s_31 + s_1614;
  assign s_31 = s_32;
  assign s_32 = s_33[23:0];
  assign s_33 = s_34 >> s_1613;
  dq #(27, 1) dq_s_34 (clk, s_34, s_35);
  assign s_35 = s_36 << s_1251;
  dq #(27, 2) dq_s_36 (clk, s_36, s_37);
  dq #(27, 1) dq_s_37 (clk, s_37, s_38);
  assign s_38 = s_39 >> s_1235;
  dq #(27, 1) dq_s_39 (clk, s_39, s_40);
  assign s_40 = s_1225?s_41:s_1223;
  assign s_41 = s_42 << s_1222;
  dq #(27, 1) dq_s_42 (clk, s_42, s_43);
  assign s_43 = s_1212?s_44:s_1210;
  assign s_44 = s_45 << s_1209;
  dq #(27, 1) dq_s_45 (clk, s_45, s_46);
  assign s_46 = s_1199?s_47:s_1197;
  assign s_47 = s_48 << s_1196;
  dq #(27, 1) dq_s_48 (clk, s_48, s_49);
  assign s_49 = s_1186?s_50:s_1184;
  assign s_50 = s_51 << s_1183;
  dq #(27, 1) dq_s_51 (clk, s_51, s_52);
  assign s_52 = s_1173?s_53:s_1171;
  assign s_53 = s_54 << s_1170;
  dq #(27, 1) dq_s_54 (clk, s_54, s_55);
  assign s_55 = s_1160?s_56:s_1158;
  assign s_56 = s_57 << s_1157;
  dq #(27, 1) dq_s_57 (clk, s_57, s_58);
  assign s_58 = s_1147?s_59:s_1145;
  assign s_59 = s_60 << s_1144;
  dq #(27, 1) dq_s_60 (clk, s_60, s_61);
  assign s_61 = s_1134?s_62:s_1132;
  assign s_62 = s_63 << s_1131;
  dq #(27, 1) dq_s_63 (clk, s_63, s_64);
  assign s_64 = s_1121?s_65:s_1119;
  assign s_65 = s_66 << s_1118;
  dq #(27, 1) dq_s_66 (clk, s_66, s_67);
  assign s_67 = s_1108?s_68:s_1106;
  assign s_68 = s_69 << s_1105;
  dq #(27, 1) dq_s_69 (clk, s_69, s_70);
  assign s_70 = s_1095?s_71:s_1093;
  assign s_71 = s_72 << s_1092;
  dq #(27, 1) dq_s_72 (clk, s_72, s_73);
  assign s_73 = s_1082?s_74:s_1080;
  assign s_74 = s_75 << s_1079;
  dq #(27, 1) dq_s_75 (clk, s_75, s_76);
  assign s_76 = s_1069?s_77:s_1067;
  assign s_77 = s_78 << s_1066;
  dq #(27, 1) dq_s_78 (clk, s_78, s_79);
  assign s_79 = s_1056?s_80:s_1054;
  assign s_80 = s_81 << s_1053;
  dq #(27, 1) dq_s_81 (clk, s_81, s_82);
  assign s_82 = s_1043?s_83:s_1041;
  assign s_83 = s_84 << s_1040;
  dq #(27, 1) dq_s_84 (clk, s_84, s_85);
  assign s_85 = s_1030?s_86:s_1028;
  assign s_86 = s_87 << s_1027;
  dq #(27, 1) dq_s_87 (clk, s_87, s_88);
  assign s_88 = s_1017?s_89:s_1015;
  assign s_89 = s_90 << s_1014;
  dq #(27, 1) dq_s_90 (clk, s_90, s_91);
  assign s_91 = s_1004?s_92:s_1002;
  assign s_92 = s_93 << s_1001;
  dq #(27, 1) dq_s_93 (clk, s_93, s_94);
  assign s_94 = s_991?s_95:s_989;
  assign s_95 = s_96 << s_988;
  dq #(27, 1) dq_s_96 (clk, s_96, s_97);
  assign s_97 = s_978?s_98:s_976;
  assign s_98 = s_99 << s_975;
  dq #(27, 1) dq_s_99 (clk, s_99, s_100);
  assign s_100 = s_965?s_101:s_963;
  assign s_101 = s_102 << s_962;
  dq #(27, 1) dq_s_102 (clk, s_102, s_103);
  assign s_103 = s_952?s_104:s_950;
  assign s_104 = s_105 << s_949;
  dq #(27, 1) dq_s_105 (clk, s_105, s_106);
  assign s_106 = s_939?s_107:s_937;
  assign s_107 = s_108 << s_936;
  dq #(27, 1) dq_s_108 (clk, s_108, s_109);
  assign s_109 = s_926?s_110:s_924;
  assign s_110 = s_111 << s_923;
  dq #(27, 1) dq_s_111 (clk, s_111, s_112);
  assign s_112 = s_913?s_113:s_911;
  assign s_113 = s_114 << s_910;
  dq #(27, 1) dq_s_114 (clk, s_114, s_115);
  assign s_115 = s_900?s_116:s_898;
  assign s_116 = s_117 << s_897;
  dq #(27, 1) dq_s_117 (clk, s_117, s_118);
  assign s_118 = s_126?s_119:s_123;
  dq #(27, 3) dq_s_119 (clk, s_119, s_120);
  assign s_120 = s_121 << s_122;
  assign s_121 = 27'd0;
  assign s_122 = 1'd1;
  dq #(27, 3) dq_s_123 (clk, s_123, s_124);
  assign s_124 = s_120 | s_125;
  assign s_125 = 1'd1;
  assign s_126 = s_127[27];
  assign s_127 = s_128 - s_513;
  assign s_128 = s_129;
  assign s_129 = s_130 << s_512;
  assign s_130 = s_131;
  dq #(24, 1) dq_s_131 (clk, s_131, s_132);
  assign s_132 = s_133 << s_144;
  dq #(24, 2) dq_s_133 (clk, s_133, s_134);
  assign s_134 = {s_135,s_143};
  assign s_135 = s_138?s_136:s_137;
  assign s_136 = 1'd0;
  assign s_137 = 1'd1;
  assign s_138 = s_139 == s_142;
  assign s_139 = s_140 - s_141;
  assign s_140 = s_5[30:23];
  assign s_141 = 7'd127;
  assign s_142 = -8'd127;
  assign s_143 = s_5[22:0];
  dq #(10, 1) dq_s_144 (clk, s_144, s_145);
  assign s_145 = s_509?s_146:s_503;
  dq #(6, 1) dq_s_146 (clk, s_146, s_147);
  assign s_147 = {s_148,s_497};
  assign s_148 = s_149 & s_331;
  assign s_149 = s_150[4];
  assign s_150 = {s_151,s_325};
  assign s_151 = s_152 & s_247;
  assign s_152 = s_153[3];
  assign s_153 = {s_154,s_241};
  assign s_154 = s_155 & s_207;
  assign s_155 = s_156[2];
  assign s_156 = {s_157,s_201};
  assign s_157 = s_158 & s_189;
  assign s_158 = s_159[1];
  assign s_159 = {s_160,s_185};
  assign s_160 = s_161 & s_183;
  assign s_161 = ~s_162;
  assign s_162 = s_163[1];
  assign s_163 = s_164[3:2];
  assign s_164 = s_165[7:4];
  assign s_165 = s_166[15:8];
  assign s_166 = s_167[31:16];
  assign s_167 = {s_168,s_182};
  assign s_168 = {s_169,s_181};
  assign s_169 = {s_170,s_180};
  assign s_170 = {s_171,s_179};
  assign s_171 = {s_172,s_178};
  assign s_172 = {s_173,s_177};
  assign s_173 = {s_174,s_176};
  assign s_174 = {s_134,s_175};
  assign s_175 = 1'd1;
  assign s_176 = 1'd1;
  assign s_177 = 1'd1;
  assign s_178 = 1'd1;
  assign s_179 = 1'd1;
  assign s_180 = 1'd1;
  assign s_181 = 1'd1;
  assign s_182 = 1'd1;
  assign s_183 = ~s_184;
  assign s_184 = s_163[0];
  assign s_185 = s_186 & s_188;
  assign s_186 = ~s_187;
  assign s_187 = s_163[1];
  assign s_188 = s_163[0];
  assign s_189 = s_190[1];
  assign s_190 = {s_191,s_197};
  assign s_191 = s_192 & s_195;
  assign s_192 = ~s_193;
  assign s_193 = s_194[1];
  assign s_194 = s_164[1:0];
  assign s_195 = ~s_196;
  assign s_196 = s_194[0];
  assign s_197 = s_198 & s_200;
  assign s_198 = ~s_199;
  assign s_199 = s_194[1];
  assign s_200 = s_194[0];
  assign s_201 = {s_202,s_204};
  assign s_202 = s_158 & s_203;
  assign s_203 = ~s_189;
  assign s_204 = s_158?s_205:s_206;
  assign s_205 = s_190[0:0];
  assign s_206 = s_159[0:0];
  assign s_207 = s_208[2];
  assign s_208 = {s_209,s_235};
  assign s_209 = s_210 & s_223;
  assign s_210 = s_211[1];
  assign s_211 = {s_212,s_219};
  assign s_212 = s_213 & s_217;
  assign s_213 = ~s_214;
  assign s_214 = s_215[1];
  assign s_215 = s_216[3:2];
  assign s_216 = s_165[3:0];
  assign s_217 = ~s_218;
  assign s_218 = s_215[0];
  assign s_219 = s_220 & s_222;
  assign s_220 = ~s_221;
  assign s_221 = s_215[1];
  assign s_222 = s_215[0];
  assign s_223 = s_224[1];
  assign s_224 = {s_225,s_231};
  assign s_225 = s_226 & s_229;
  assign s_226 = ~s_227;
  assign s_227 = s_228[1];
  assign s_228 = s_216[1:0];
  assign s_229 = ~s_230;
  assign s_230 = s_228[0];
  assign s_231 = s_232 & s_234;
  assign s_232 = ~s_233;
  assign s_233 = s_228[1];
  assign s_234 = s_228[0];
  assign s_235 = {s_236,s_238};
  assign s_236 = s_210 & s_237;
  assign s_237 = ~s_223;
  assign s_238 = s_210?s_239:s_240;
  assign s_239 = s_224[0:0];
  assign s_240 = s_211[0:0];
  assign s_241 = {s_242,s_244};
  assign s_242 = s_155 & s_243;
  assign s_243 = ~s_207;
  assign s_244 = s_155?s_245:s_246;
  assign s_245 = s_208[1:0];
  assign s_246 = s_156[1:0];
  assign s_247 = s_248[3];
  assign s_248 = {s_249,s_319};
  assign s_249 = s_250 & s_285;
  assign s_250 = s_251[2];
  assign s_251 = {s_252,s_279};
  assign s_252 = s_253 & s_267;
  assign s_253 = s_254[1];
  assign s_254 = {s_255,s_263};
  assign s_255 = s_256 & s_261;
  assign s_256 = ~s_257;
  assign s_257 = s_258[1];
  assign s_258 = s_259[3:2];
  assign s_259 = s_260[7:4];
  assign s_260 = s_166[7:0];
  assign s_261 = ~s_262;
  assign s_262 = s_258[0];
  assign s_263 = s_264 & s_266;
  assign s_264 = ~s_265;
  assign s_265 = s_258[1];
  assign s_266 = s_258[0];
  assign s_267 = s_268[1];
  assign s_268 = {s_269,s_275};
  assign s_269 = s_270 & s_273;
  assign s_270 = ~s_271;
  assign s_271 = s_272[1];
  assign s_272 = s_259[1:0];
  assign s_273 = ~s_274;
  assign s_274 = s_272[0];
  assign s_275 = s_276 & s_278;
  assign s_276 = ~s_277;
  assign s_277 = s_272[1];
  assign s_278 = s_272[0];
  assign s_279 = {s_280,s_282};
  assign s_280 = s_253 & s_281;
  assign s_281 = ~s_267;
  assign s_282 = s_253?s_283:s_284;
  assign s_283 = s_268[0:0];
  assign s_284 = s_254[0:0];
  assign s_285 = s_286[2];
  assign s_286 = {s_287,s_313};
  assign s_287 = s_288 & s_301;
  assign s_288 = s_289[1];
  assign s_289 = {s_290,s_297};
  assign s_290 = s_291 & s_295;
  assign s_291 = ~s_292;
  assign s_292 = s_293[1];
  assign s_293 = s_294[3:2];
  assign s_294 = s_260[3:0];
  assign s_295 = ~s_296;
  assign s_296 = s_293[0];
  assign s_297 = s_298 & s_300;
  assign s_298 = ~s_299;
  assign s_299 = s_293[1];
  assign s_300 = s_293[0];
  assign s_301 = s_302[1];
  assign s_302 = {s_303,s_309};
  assign s_303 = s_304 & s_307;
  assign s_304 = ~s_305;
  assign s_305 = s_306[1];
  assign s_306 = s_294[1:0];
  assign s_307 = ~s_308;
  assign s_308 = s_306[0];
  assign s_309 = s_310 & s_312;
  assign s_310 = ~s_311;
  assign s_311 = s_306[1];
  assign s_312 = s_306[0];
  assign s_313 = {s_314,s_316};
  assign s_314 = s_288 & s_315;
  assign s_315 = ~s_301;
  assign s_316 = s_288?s_317:s_318;
  assign s_317 = s_302[0:0];
  assign s_318 = s_289[0:0];
  assign s_319 = {s_320,s_322};
  assign s_320 = s_250 & s_321;
  assign s_321 = ~s_285;
  assign s_322 = s_250?s_323:s_324;
  assign s_323 = s_286[1:0];
  assign s_324 = s_251[1:0];
  assign s_325 = {s_326,s_328};
  assign s_326 = s_152 & s_327;
  assign s_327 = ~s_247;
  assign s_328 = s_152?s_329:s_330;
  assign s_329 = s_248[2:0];
  assign s_330 = s_153[2:0];
  assign s_331 = s_332[4];
  assign s_332 = {s_333,s_491};
  assign s_333 = s_334 & s_413;
  assign s_334 = s_335[3];
  assign s_335 = {s_336,s_407};
  assign s_336 = s_337 & s_373;
  assign s_337 = s_338[2];
  assign s_338 = {s_339,s_367};
  assign s_339 = s_340 & s_355;
  assign s_340 = s_341[1];
  assign s_341 = {s_342,s_351};
  assign s_342 = s_343 & s_349;
  assign s_343 = ~s_344;
  assign s_344 = s_345[1];
  assign s_345 = s_346[3:2];
  assign s_346 = s_347[7:4];
  assign s_347 = s_348[15:8];
  assign s_348 = s_167[15:0];
  assign s_349 = ~s_350;
  assign s_350 = s_345[0];
  assign s_351 = s_352 & s_354;
  assign s_352 = ~s_353;
  assign s_353 = s_345[1];
  assign s_354 = s_345[0];
  assign s_355 = s_356[1];
  assign s_356 = {s_357,s_363};
  assign s_357 = s_358 & s_361;
  assign s_358 = ~s_359;
  assign s_359 = s_360[1];
  assign s_360 = s_346[1:0];
  assign s_361 = ~s_362;
  assign s_362 = s_360[0];
  assign s_363 = s_364 & s_366;
  assign s_364 = ~s_365;
  assign s_365 = s_360[1];
  assign s_366 = s_360[0];
  assign s_367 = {s_368,s_370};
  assign s_368 = s_340 & s_369;
  assign s_369 = ~s_355;
  assign s_370 = s_340?s_371:s_372;
  assign s_371 = s_356[0:0];
  assign s_372 = s_341[0:0];
  assign s_373 = s_374[2];
  assign s_374 = {s_375,s_401};
  assign s_375 = s_376 & s_389;
  assign s_376 = s_377[1];
  assign s_377 = {s_378,s_385};
  assign s_378 = s_379 & s_383;
  assign s_379 = ~s_380;
  assign s_380 = s_381[1];
  assign s_381 = s_382[3:2];
  assign s_382 = s_347[3:0];
  assign s_383 = ~s_384;
  assign s_384 = s_381[0];
  assign s_385 = s_386 & s_388;
  assign s_386 = ~s_387;
  assign s_387 = s_381[1];
  assign s_388 = s_381[0];
  assign s_389 = s_390[1];
  assign s_390 = {s_391,s_397};
  assign s_391 = s_392 & s_395;
  assign s_392 = ~s_393;
  assign s_393 = s_394[1];
  assign s_394 = s_382[1:0];
  assign s_395 = ~s_396;
  assign s_396 = s_394[0];
  assign s_397 = s_398 & s_400;
  assign s_398 = ~s_399;
  assign s_399 = s_394[1];
  assign s_400 = s_394[0];
  assign s_401 = {s_402,s_404};
  assign s_402 = s_376 & s_403;
  assign s_403 = ~s_389;
  assign s_404 = s_376?s_405:s_406;
  assign s_405 = s_390[0:0];
  assign s_406 = s_377[0:0];
  assign s_407 = {s_408,s_410};
  assign s_408 = s_337 & s_409;
  assign s_409 = ~s_373;
  assign s_410 = s_337?s_411:s_412;
  assign s_411 = s_374[1:0];
  assign s_412 = s_338[1:0];
  assign s_413 = s_414[3];
  assign s_414 = {s_415,s_485};
  assign s_415 = s_416 & s_451;
  assign s_416 = s_417[2];
  assign s_417 = {s_418,s_445};
  assign s_418 = s_419 & s_433;
  assign s_419 = s_420[1];
  assign s_420 = {s_421,s_429};
  assign s_421 = s_422 & s_427;
  assign s_422 = ~s_423;
  assign s_423 = s_424[1];
  assign s_424 = s_425[3:2];
  assign s_425 = s_426[7:4];
  assign s_426 = s_348[7:0];
  assign s_427 = ~s_428;
  assign s_428 = s_424[0];
  assign s_429 = s_430 & s_432;
  assign s_430 = ~s_431;
  assign s_431 = s_424[1];
  assign s_432 = s_424[0];
  assign s_433 = s_434[1];
  assign s_434 = {s_435,s_441};
  assign s_435 = s_436 & s_439;
  assign s_436 = ~s_437;
  assign s_437 = s_438[1];
  assign s_438 = s_425[1:0];
  assign s_439 = ~s_440;
  assign s_440 = s_438[0];
  assign s_441 = s_442 & s_444;
  assign s_442 = ~s_443;
  assign s_443 = s_438[1];
  assign s_444 = s_438[0];
  assign s_445 = {s_446,s_448};
  assign s_446 = s_419 & s_447;
  assign s_447 = ~s_433;
  assign s_448 = s_419?s_449:s_450;
  assign s_449 = s_434[0:0];
  assign s_450 = s_420[0:0];
  assign s_451 = s_452[2];
  assign s_452 = {s_453,s_479};
  assign s_453 = s_454 & s_467;
  assign s_454 = s_455[1];
  assign s_455 = {s_456,s_463};
  assign s_456 = s_457 & s_461;
  assign s_457 = ~s_458;
  assign s_458 = s_459[1];
  assign s_459 = s_460[3:2];
  assign s_460 = s_426[3:0];
  assign s_461 = ~s_462;
  assign s_462 = s_459[0];
  assign s_463 = s_464 & s_466;
  assign s_464 = ~s_465;
  assign s_465 = s_459[1];
  assign s_466 = s_459[0];
  assign s_467 = s_468[1];
  assign s_468 = {s_469,s_475};
  assign s_469 = s_470 & s_473;
  assign s_470 = ~s_471;
  assign s_471 = s_472[1];
  assign s_472 = s_460[1:0];
  assign s_473 = ~s_474;
  assign s_474 = s_472[0];
  assign s_475 = s_476 & s_478;
  assign s_476 = ~s_477;
  assign s_477 = s_472[1];
  assign s_478 = s_472[0];
  assign s_479 = {s_480,s_482};
  assign s_480 = s_454 & s_481;
  assign s_481 = ~s_467;
  assign s_482 = s_454?s_483:s_484;
  assign s_483 = s_468[0:0];
  assign s_484 = s_455[0:0];
  assign s_485 = {s_486,s_488};
  assign s_486 = s_416 & s_487;
  assign s_487 = ~s_451;
  assign s_488 = s_416?s_489:s_490;
  assign s_489 = s_452[1:0];
  assign s_490 = s_417[1:0];
  assign s_491 = {s_492,s_494};
  assign s_492 = s_334 & s_493;
  assign s_493 = ~s_413;
  assign s_494 = s_334?s_495:s_496;
  assign s_495 = s_414[2:0];
  assign s_496 = s_335[2:0];
  assign s_497 = {s_498,s_500};
  assign s_498 = s_149 & s_499;
  assign s_499 = ~s_331;
  assign s_500 = s_149?s_501:s_502;
  assign s_501 = s_332[3:0];
  assign s_502 = s_150[3:0];
  dq #(10, 1) dq_s_503 (clk, s_503, s_504);
  assign s_504 = s_505 - s_508;
  assign s_505 = $signed(s_506);
  assign s_506 = s_138?s_507:s_139;
  assign s_507 = -8'd126;
  assign s_508 = -10'd252;
  assign s_509 = s_510 <= s_511;
  assign s_510 = s_146;
  dq #(10, 1) dq_s_511 (clk, s_511, s_504);
  assign s_512 = 2'd3;
  assign s_513 = s_514 << s_896;
  assign s_514 = s_515;
  dq #(24, 1) dq_s_515 (clk, s_515, s_516);
  assign s_516 = s_517 << s_528;
  dq #(24, 2) dq_s_517 (clk, s_517, s_518);
  assign s_518 = {s_519,s_527};
  assign s_519 = s_522?s_520:s_521;
  assign s_520 = 1'd0;
  assign s_521 = 1'd1;
  assign s_522 = s_523 == s_526;
  assign s_523 = s_524 - s_525;
  assign s_524 = s_7[30:23];
  assign s_525 = 7'd127;
  assign s_526 = -8'd127;
  assign s_527 = s_7[22:0];
  dq #(10, 1) dq_s_528 (clk, s_528, s_529);
  assign s_529 = s_893?s_530:s_887;
  dq #(6, 1) dq_s_530 (clk, s_530, s_531);
  assign s_531 = {s_532,s_881};
  assign s_532 = s_533 & s_715;
  assign s_533 = s_534[4];
  assign s_534 = {s_535,s_709};
  assign s_535 = s_536 & s_631;
  assign s_536 = s_537[3];
  assign s_537 = {s_538,s_625};
  assign s_538 = s_539 & s_591;
  assign s_539 = s_540[2];
  assign s_540 = {s_541,s_585};
  assign s_541 = s_542 & s_573;
  assign s_542 = s_543[1];
  assign s_543 = {s_544,s_569};
  assign s_544 = s_545 & s_567;
  assign s_545 = ~s_546;
  assign s_546 = s_547[1];
  assign s_547 = s_548[3:2];
  assign s_548 = s_549[7:4];
  assign s_549 = s_550[15:8];
  assign s_550 = s_551[31:16];
  assign s_551 = {s_552,s_566};
  assign s_552 = {s_553,s_565};
  assign s_553 = {s_554,s_564};
  assign s_554 = {s_555,s_563};
  assign s_555 = {s_556,s_562};
  assign s_556 = {s_557,s_561};
  assign s_557 = {s_558,s_560};
  assign s_558 = {s_518,s_559};
  assign s_559 = 1'd1;
  assign s_560 = 1'd1;
  assign s_561 = 1'd1;
  assign s_562 = 1'd1;
  assign s_563 = 1'd1;
  assign s_564 = 1'd1;
  assign s_565 = 1'd1;
  assign s_566 = 1'd1;
  assign s_567 = ~s_568;
  assign s_568 = s_547[0];
  assign s_569 = s_570 & s_572;
  assign s_570 = ~s_571;
  assign s_571 = s_547[1];
  assign s_572 = s_547[0];
  assign s_573 = s_574[1];
  assign s_574 = {s_575,s_581};
  assign s_575 = s_576 & s_579;
  assign s_576 = ~s_577;
  assign s_577 = s_578[1];
  assign s_578 = s_548[1:0];
  assign s_579 = ~s_580;
  assign s_580 = s_578[0];
  assign s_581 = s_582 & s_584;
  assign s_582 = ~s_583;
  assign s_583 = s_578[1];
  assign s_584 = s_578[0];
  assign s_585 = {s_586,s_588};
  assign s_586 = s_542 & s_587;
  assign s_587 = ~s_573;
  assign s_588 = s_542?s_589:s_590;
  assign s_589 = s_574[0:0];
  assign s_590 = s_543[0:0];
  assign s_591 = s_592[2];
  assign s_592 = {s_593,s_619};
  assign s_593 = s_594 & s_607;
  assign s_594 = s_595[1];
  assign s_595 = {s_596,s_603};
  assign s_596 = s_597 & s_601;
  assign s_597 = ~s_598;
  assign s_598 = s_599[1];
  assign s_599 = s_600[3:2];
  assign s_600 = s_549[3:0];
  assign s_601 = ~s_602;
  assign s_602 = s_599[0];
  assign s_603 = s_604 & s_606;
  assign s_604 = ~s_605;
  assign s_605 = s_599[1];
  assign s_606 = s_599[0];
  assign s_607 = s_608[1];
  assign s_608 = {s_609,s_615};
  assign s_609 = s_610 & s_613;
  assign s_610 = ~s_611;
  assign s_611 = s_612[1];
  assign s_612 = s_600[1:0];
  assign s_613 = ~s_614;
  assign s_614 = s_612[0];
  assign s_615 = s_616 & s_618;
  assign s_616 = ~s_617;
  assign s_617 = s_612[1];
  assign s_618 = s_612[0];
  assign s_619 = {s_620,s_622};
  assign s_620 = s_594 & s_621;
  assign s_621 = ~s_607;
  assign s_622 = s_594?s_623:s_624;
  assign s_623 = s_608[0:0];
  assign s_624 = s_595[0:0];
  assign s_625 = {s_626,s_628};
  assign s_626 = s_539 & s_627;
  assign s_627 = ~s_591;
  assign s_628 = s_539?s_629:s_630;
  assign s_629 = s_592[1:0];
  assign s_630 = s_540[1:0];
  assign s_631 = s_632[3];
  assign s_632 = {s_633,s_703};
  assign s_633 = s_634 & s_669;
  assign s_634 = s_635[2];
  assign s_635 = {s_636,s_663};
  assign s_636 = s_637 & s_651;
  assign s_637 = s_638[1];
  assign s_638 = {s_639,s_647};
  assign s_639 = s_640 & s_645;
  assign s_640 = ~s_641;
  assign s_641 = s_642[1];
  assign s_642 = s_643[3:2];
  assign s_643 = s_644[7:4];
  assign s_644 = s_550[7:0];
  assign s_645 = ~s_646;
  assign s_646 = s_642[0];
  assign s_647 = s_648 & s_650;
  assign s_648 = ~s_649;
  assign s_649 = s_642[1];
  assign s_650 = s_642[0];
  assign s_651 = s_652[1];
  assign s_652 = {s_653,s_659};
  assign s_653 = s_654 & s_657;
  assign s_654 = ~s_655;
  assign s_655 = s_656[1];
  assign s_656 = s_643[1:0];
  assign s_657 = ~s_658;
  assign s_658 = s_656[0];
  assign s_659 = s_660 & s_662;
  assign s_660 = ~s_661;
  assign s_661 = s_656[1];
  assign s_662 = s_656[0];
  assign s_663 = {s_664,s_666};
  assign s_664 = s_637 & s_665;
  assign s_665 = ~s_651;
  assign s_666 = s_637?s_667:s_668;
  assign s_667 = s_652[0:0];
  assign s_668 = s_638[0:0];
  assign s_669 = s_670[2];
  assign s_670 = {s_671,s_697};
  assign s_671 = s_672 & s_685;
  assign s_672 = s_673[1];
  assign s_673 = {s_674,s_681};
  assign s_674 = s_675 & s_679;
  assign s_675 = ~s_676;
  assign s_676 = s_677[1];
  assign s_677 = s_678[3:2];
  assign s_678 = s_644[3:0];
  assign s_679 = ~s_680;
  assign s_680 = s_677[0];
  assign s_681 = s_682 & s_684;
  assign s_682 = ~s_683;
  assign s_683 = s_677[1];
  assign s_684 = s_677[0];
  assign s_685 = s_686[1];
  assign s_686 = {s_687,s_693};
  assign s_687 = s_688 & s_691;
  assign s_688 = ~s_689;
  assign s_689 = s_690[1];
  assign s_690 = s_678[1:0];
  assign s_691 = ~s_692;
  assign s_692 = s_690[0];
  assign s_693 = s_694 & s_696;
  assign s_694 = ~s_695;
  assign s_695 = s_690[1];
  assign s_696 = s_690[0];
  assign s_697 = {s_698,s_700};
  assign s_698 = s_672 & s_699;
  assign s_699 = ~s_685;
  assign s_700 = s_672?s_701:s_702;
  assign s_701 = s_686[0:0];
  assign s_702 = s_673[0:0];
  assign s_703 = {s_704,s_706};
  assign s_704 = s_634 & s_705;
  assign s_705 = ~s_669;
  assign s_706 = s_634?s_707:s_708;
  assign s_707 = s_670[1:0];
  assign s_708 = s_635[1:0];
  assign s_709 = {s_710,s_712};
  assign s_710 = s_536 & s_711;
  assign s_711 = ~s_631;
  assign s_712 = s_536?s_713:s_714;
  assign s_713 = s_632[2:0];
  assign s_714 = s_537[2:0];
  assign s_715 = s_716[4];
  assign s_716 = {s_717,s_875};
  assign s_717 = s_718 & s_797;
  assign s_718 = s_719[3];
  assign s_719 = {s_720,s_791};
  assign s_720 = s_721 & s_757;
  assign s_721 = s_722[2];
  assign s_722 = {s_723,s_751};
  assign s_723 = s_724 & s_739;
  assign s_724 = s_725[1];
  assign s_725 = {s_726,s_735};
  assign s_726 = s_727 & s_733;
  assign s_727 = ~s_728;
  assign s_728 = s_729[1];
  assign s_729 = s_730[3:2];
  assign s_730 = s_731[7:4];
  assign s_731 = s_732[15:8];
  assign s_732 = s_551[15:0];
  assign s_733 = ~s_734;
  assign s_734 = s_729[0];
  assign s_735 = s_736 & s_738;
  assign s_736 = ~s_737;
  assign s_737 = s_729[1];
  assign s_738 = s_729[0];
  assign s_739 = s_740[1];
  assign s_740 = {s_741,s_747};
  assign s_741 = s_742 & s_745;
  assign s_742 = ~s_743;
  assign s_743 = s_744[1];
  assign s_744 = s_730[1:0];
  assign s_745 = ~s_746;
  assign s_746 = s_744[0];
  assign s_747 = s_748 & s_750;
  assign s_748 = ~s_749;
  assign s_749 = s_744[1];
  assign s_750 = s_744[0];
  assign s_751 = {s_752,s_754};
  assign s_752 = s_724 & s_753;
  assign s_753 = ~s_739;
  assign s_754 = s_724?s_755:s_756;
  assign s_755 = s_740[0:0];
  assign s_756 = s_725[0:0];
  assign s_757 = s_758[2];
  assign s_758 = {s_759,s_785};
  assign s_759 = s_760 & s_773;
  assign s_760 = s_761[1];
  assign s_761 = {s_762,s_769};
  assign s_762 = s_763 & s_767;
  assign s_763 = ~s_764;
  assign s_764 = s_765[1];
  assign s_765 = s_766[3:2];
  assign s_766 = s_731[3:0];
  assign s_767 = ~s_768;
  assign s_768 = s_765[0];
  assign s_769 = s_770 & s_772;
  assign s_770 = ~s_771;
  assign s_771 = s_765[1];
  assign s_772 = s_765[0];
  assign s_773 = s_774[1];
  assign s_774 = {s_775,s_781};
  assign s_775 = s_776 & s_779;
  assign s_776 = ~s_777;
  assign s_777 = s_778[1];
  assign s_778 = s_766[1:0];
  assign s_779 = ~s_780;
  assign s_780 = s_778[0];
  assign s_781 = s_782 & s_784;
  assign s_782 = ~s_783;
  assign s_783 = s_778[1];
  assign s_784 = s_778[0];
  assign s_785 = {s_786,s_788};
  assign s_786 = s_760 & s_787;
  assign s_787 = ~s_773;
  assign s_788 = s_760?s_789:s_790;
  assign s_789 = s_774[0:0];
  assign s_790 = s_761[0:0];
  assign s_791 = {s_792,s_794};
  assign s_792 = s_721 & s_793;
  assign s_793 = ~s_757;
  assign s_794 = s_721?s_795:s_796;
  assign s_795 = s_758[1:0];
  assign s_796 = s_722[1:0];
  assign s_797 = s_798[3];
  assign s_798 = {s_799,s_869};
  assign s_799 = s_800 & s_835;
  assign s_800 = s_801[2];
  assign s_801 = {s_802,s_829};
  assign s_802 = s_803 & s_817;
  assign s_803 = s_804[1];
  assign s_804 = {s_805,s_813};
  assign s_805 = s_806 & s_811;
  assign s_806 = ~s_807;
  assign s_807 = s_808[1];
  assign s_808 = s_809[3:2];
  assign s_809 = s_810[7:4];
  assign s_810 = s_732[7:0];
  assign s_811 = ~s_812;
  assign s_812 = s_808[0];
  assign s_813 = s_814 & s_816;
  assign s_814 = ~s_815;
  assign s_815 = s_808[1];
  assign s_816 = s_808[0];
  assign s_817 = s_818[1];
  assign s_818 = {s_819,s_825};
  assign s_819 = s_820 & s_823;
  assign s_820 = ~s_821;
  assign s_821 = s_822[1];
  assign s_822 = s_809[1:0];
  assign s_823 = ~s_824;
  assign s_824 = s_822[0];
  assign s_825 = s_826 & s_828;
  assign s_826 = ~s_827;
  assign s_827 = s_822[1];
  assign s_828 = s_822[0];
  assign s_829 = {s_830,s_832};
  assign s_830 = s_803 & s_831;
  assign s_831 = ~s_817;
  assign s_832 = s_803?s_833:s_834;
  assign s_833 = s_818[0:0];
  assign s_834 = s_804[0:0];
  assign s_835 = s_836[2];
  assign s_836 = {s_837,s_863};
  assign s_837 = s_838 & s_851;
  assign s_838 = s_839[1];
  assign s_839 = {s_840,s_847};
  assign s_840 = s_841 & s_845;
  assign s_841 = ~s_842;
  assign s_842 = s_843[1];
  assign s_843 = s_844[3:2];
  assign s_844 = s_810[3:0];
  assign s_845 = ~s_846;
  assign s_846 = s_843[0];
  assign s_847 = s_848 & s_850;
  assign s_848 = ~s_849;
  assign s_849 = s_843[1];
  assign s_850 = s_843[0];
  assign s_851 = s_852[1];
  assign s_852 = {s_853,s_859};
  assign s_853 = s_854 & s_857;
  assign s_854 = ~s_855;
  assign s_855 = s_856[1];
  assign s_856 = s_844[1:0];
  assign s_857 = ~s_858;
  assign s_858 = s_856[0];
  assign s_859 = s_860 & s_862;
  assign s_860 = ~s_861;
  assign s_861 = s_856[1];
  assign s_862 = s_856[0];
  assign s_863 = {s_864,s_866};
  assign s_864 = s_838 & s_865;
  assign s_865 = ~s_851;
  assign s_866 = s_838?s_867:s_868;
  assign s_867 = s_852[0:0];
  assign s_868 = s_839[0:0];
  assign s_869 = {s_870,s_872};
  assign s_870 = s_800 & s_871;
  assign s_871 = ~s_835;
  assign s_872 = s_800?s_873:s_874;
  assign s_873 = s_836[1:0];
  assign s_874 = s_801[1:0];
  assign s_875 = {s_876,s_878};
  assign s_876 = s_718 & s_877;
  assign s_877 = ~s_797;
  assign s_878 = s_718?s_879:s_880;
  assign s_879 = s_798[2:0];
  assign s_880 = s_719[2:0];
  assign s_881 = {s_882,s_884};
  assign s_882 = s_533 & s_883;
  assign s_883 = ~s_715;
  assign s_884 = s_533?s_885:s_886;
  assign s_885 = s_716[3:0];
  assign s_886 = s_534[3:0];
  dq #(10, 1) dq_s_887 (clk, s_887, s_888);
  assign s_888 = s_889 - s_892;
  assign s_889 = $signed(s_890);
  assign s_890 = s_522?s_891:s_523;
  assign s_891 = -8'd126;
  assign s_892 = -10'd252;
  assign s_893 = s_894 <= s_895;
  assign s_894 = s_530;
  dq #(10, 1) dq_s_895 (clk, s_895, s_888);
  assign s_896 = 2'd3;
  assign s_897 = 1'd1;
  assign s_898 = s_116 | s_899;
  assign s_899 = 1'd1;
  assign s_900 = s_901[27];
  assign s_901 = s_902 - s_909;
  assign s_902 = s_903;
  assign s_903 = s_904 | s_908;
  assign s_904 = s_905 << s_907;
  dq #(28, 1) dq_s_905 (clk, s_905, s_906);
  assign s_906 = s_126?s_129:s_127;
  assign s_907 = 1'd1;
  assign s_908 = 1'd0;
  dq #(27, 1) dq_s_909 (clk, s_909, s_513);
  assign s_910 = 1'd1;
  assign s_911 = s_113 | s_912;
  assign s_912 = 1'd1;
  assign s_913 = s_914[27];
  assign s_914 = s_915 - s_922;
  assign s_915 = s_916;
  assign s_916 = s_917 | s_921;
  assign s_917 = s_918 << s_920;
  dq #(28, 1) dq_s_918 (clk, s_918, s_919);
  assign s_919 = s_900?s_903:s_901;
  assign s_920 = 1'd1;
  assign s_921 = 1'd0;
  dq #(27, 2) dq_s_922 (clk, s_922, s_513);
  assign s_923 = 1'd1;
  assign s_924 = s_110 | s_925;
  assign s_925 = 1'd1;
  assign s_926 = s_927[27];
  assign s_927 = s_928 - s_935;
  assign s_928 = s_929;
  assign s_929 = s_930 | s_934;
  assign s_930 = s_931 << s_933;
  dq #(28, 1) dq_s_931 (clk, s_931, s_932);
  assign s_932 = s_913?s_916:s_914;
  assign s_933 = 1'd1;
  assign s_934 = 1'd0;
  dq #(27, 3) dq_s_935 (clk, s_935, s_513);
  assign s_936 = 1'd1;
  assign s_937 = s_107 | s_938;
  assign s_938 = 1'd1;
  assign s_939 = s_940[27];
  assign s_940 = s_941 - s_948;
  assign s_941 = s_942;
  assign s_942 = s_943 | s_947;
  assign s_943 = s_944 << s_946;
  dq #(28, 1) dq_s_944 (clk, s_944, s_945);
  assign s_945 = s_926?s_929:s_927;
  assign s_946 = 1'd1;
  assign s_947 = 1'd0;
  dq #(27, 4) dq_s_948 (clk, s_948, s_513);
  assign s_949 = 1'd1;
  assign s_950 = s_104 | s_951;
  assign s_951 = 1'd1;
  assign s_952 = s_953[27];
  assign s_953 = s_954 - s_961;
  assign s_954 = s_955;
  assign s_955 = s_956 | s_960;
  assign s_956 = s_957 << s_959;
  dq #(28, 1) dq_s_957 (clk, s_957, s_958);
  assign s_958 = s_939?s_942:s_940;
  assign s_959 = 1'd1;
  assign s_960 = 1'd0;
  dq #(27, 5) dq_s_961 (clk, s_961, s_513);
  assign s_962 = 1'd1;
  assign s_963 = s_101 | s_964;
  assign s_964 = 1'd1;
  assign s_965 = s_966[27];
  assign s_966 = s_967 - s_974;
  assign s_967 = s_968;
  assign s_968 = s_969 | s_973;
  assign s_969 = s_970 << s_972;
  dq #(28, 1) dq_s_970 (clk, s_970, s_971);
  assign s_971 = s_952?s_955:s_953;
  assign s_972 = 1'd1;
  assign s_973 = 1'd0;
  dq #(27, 6) dq_s_974 (clk, s_974, s_513);
  assign s_975 = 1'd1;
  assign s_976 = s_98 | s_977;
  assign s_977 = 1'd1;
  assign s_978 = s_979[27];
  assign s_979 = s_980 - s_987;
  assign s_980 = s_981;
  assign s_981 = s_982 | s_986;
  assign s_982 = s_983 << s_985;
  dq #(28, 1) dq_s_983 (clk, s_983, s_984);
  assign s_984 = s_965?s_968:s_966;
  assign s_985 = 1'd1;
  assign s_986 = 1'd0;
  dq #(27, 7) dq_s_987 (clk, s_987, s_513);
  assign s_988 = 1'd1;
  assign s_989 = s_95 | s_990;
  assign s_990 = 1'd1;
  assign s_991 = s_992[27];
  assign s_992 = s_993 - s_1000;
  assign s_993 = s_994;
  assign s_994 = s_995 | s_999;
  assign s_995 = s_996 << s_998;
  dq #(28, 1) dq_s_996 (clk, s_996, s_997);
  assign s_997 = s_978?s_981:s_979;
  assign s_998 = 1'd1;
  assign s_999 = 1'd0;
  dq #(27, 8) dq_s_1000 (clk, s_1000, s_513);
  assign s_1001 = 1'd1;
  assign s_1002 = s_92 | s_1003;
  assign s_1003 = 1'd1;
  assign s_1004 = s_1005[27];
  assign s_1005 = s_1006 - s_1013;
  assign s_1006 = s_1007;
  assign s_1007 = s_1008 | s_1012;
  assign s_1008 = s_1009 << s_1011;
  dq #(28, 1) dq_s_1009 (clk, s_1009, s_1010);
  assign s_1010 = s_991?s_994:s_992;
  assign s_1011 = 1'd1;
  assign s_1012 = 1'd0;
  dq #(27, 9) dq_s_1013 (clk, s_1013, s_513);
  assign s_1014 = 1'd1;
  assign s_1015 = s_89 | s_1016;
  assign s_1016 = 1'd1;
  assign s_1017 = s_1018[27];
  assign s_1018 = s_1019 - s_1026;
  assign s_1019 = s_1020;
  assign s_1020 = s_1021 | s_1025;
  assign s_1021 = s_1022 << s_1024;
  dq #(28, 1) dq_s_1022 (clk, s_1022, s_1023);
  assign s_1023 = s_1004?s_1007:s_1005;
  assign s_1024 = 1'd1;
  assign s_1025 = 1'd0;
  dq #(27, 10) dq_s_1026 (clk, s_1026, s_513);
  assign s_1027 = 1'd1;
  assign s_1028 = s_86 | s_1029;
  assign s_1029 = 1'd1;
  assign s_1030 = s_1031[27];
  assign s_1031 = s_1032 - s_1039;
  assign s_1032 = s_1033;
  assign s_1033 = s_1034 | s_1038;
  assign s_1034 = s_1035 << s_1037;
  dq #(28, 1) dq_s_1035 (clk, s_1035, s_1036);
  assign s_1036 = s_1017?s_1020:s_1018;
  assign s_1037 = 1'd1;
  assign s_1038 = 1'd0;
  dq #(27, 11) dq_s_1039 (clk, s_1039, s_513);
  assign s_1040 = 1'd1;
  assign s_1041 = s_83 | s_1042;
  assign s_1042 = 1'd1;
  assign s_1043 = s_1044[27];
  assign s_1044 = s_1045 - s_1052;
  assign s_1045 = s_1046;
  assign s_1046 = s_1047 | s_1051;
  assign s_1047 = s_1048 << s_1050;
  dq #(28, 1) dq_s_1048 (clk, s_1048, s_1049);
  assign s_1049 = s_1030?s_1033:s_1031;
  assign s_1050 = 1'd1;
  assign s_1051 = 1'd0;
  dq #(27, 12) dq_s_1052 (clk, s_1052, s_513);
  assign s_1053 = 1'd1;
  assign s_1054 = s_80 | s_1055;
  assign s_1055 = 1'd1;
  assign s_1056 = s_1057[27];
  assign s_1057 = s_1058 - s_1065;
  assign s_1058 = s_1059;
  assign s_1059 = s_1060 | s_1064;
  assign s_1060 = s_1061 << s_1063;
  dq #(28, 1) dq_s_1061 (clk, s_1061, s_1062);
  assign s_1062 = s_1043?s_1046:s_1044;
  assign s_1063 = 1'd1;
  assign s_1064 = 1'd0;
  dq #(27, 13) dq_s_1065 (clk, s_1065, s_513);
  assign s_1066 = 1'd1;
  assign s_1067 = s_77 | s_1068;
  assign s_1068 = 1'd1;
  assign s_1069 = s_1070[27];
  assign s_1070 = s_1071 - s_1078;
  assign s_1071 = s_1072;
  assign s_1072 = s_1073 | s_1077;
  assign s_1073 = s_1074 << s_1076;
  dq #(28, 1) dq_s_1074 (clk, s_1074, s_1075);
  assign s_1075 = s_1056?s_1059:s_1057;
  assign s_1076 = 1'd1;
  assign s_1077 = 1'd0;
  dq #(27, 14) dq_s_1078 (clk, s_1078, s_513);
  assign s_1079 = 1'd1;
  assign s_1080 = s_74 | s_1081;
  assign s_1081 = 1'd1;
  assign s_1082 = s_1083[27];
  assign s_1083 = s_1084 - s_1091;
  assign s_1084 = s_1085;
  assign s_1085 = s_1086 | s_1090;
  assign s_1086 = s_1087 << s_1089;
  dq #(28, 1) dq_s_1087 (clk, s_1087, s_1088);
  assign s_1088 = s_1069?s_1072:s_1070;
  assign s_1089 = 1'd1;
  assign s_1090 = 1'd0;
  dq #(27, 15) dq_s_1091 (clk, s_1091, s_513);
  assign s_1092 = 1'd1;
  assign s_1093 = s_71 | s_1094;
  assign s_1094 = 1'd1;
  assign s_1095 = s_1096[27];
  assign s_1096 = s_1097 - s_1104;
  assign s_1097 = s_1098;
  assign s_1098 = s_1099 | s_1103;
  assign s_1099 = s_1100 << s_1102;
  dq #(28, 1) dq_s_1100 (clk, s_1100, s_1101);
  assign s_1101 = s_1082?s_1085:s_1083;
  assign s_1102 = 1'd1;
  assign s_1103 = 1'd0;
  dq #(27, 16) dq_s_1104 (clk, s_1104, s_513);
  assign s_1105 = 1'd1;
  assign s_1106 = s_68 | s_1107;
  assign s_1107 = 1'd1;
  assign s_1108 = s_1109[27];
  assign s_1109 = s_1110 - s_1117;
  assign s_1110 = s_1111;
  assign s_1111 = s_1112 | s_1116;
  assign s_1112 = s_1113 << s_1115;
  dq #(28, 1) dq_s_1113 (clk, s_1113, s_1114);
  assign s_1114 = s_1095?s_1098:s_1096;
  assign s_1115 = 1'd1;
  assign s_1116 = 1'd0;
  dq #(27, 17) dq_s_1117 (clk, s_1117, s_513);
  assign s_1118 = 1'd1;
  assign s_1119 = s_65 | s_1120;
  assign s_1120 = 1'd1;
  assign s_1121 = s_1122[27];
  assign s_1122 = s_1123 - s_1130;
  assign s_1123 = s_1124;
  assign s_1124 = s_1125 | s_1129;
  assign s_1125 = s_1126 << s_1128;
  dq #(28, 1) dq_s_1126 (clk, s_1126, s_1127);
  assign s_1127 = s_1108?s_1111:s_1109;
  assign s_1128 = 1'd1;
  assign s_1129 = 1'd0;
  dq #(27, 18) dq_s_1130 (clk, s_1130, s_513);
  assign s_1131 = 1'd1;
  assign s_1132 = s_62 | s_1133;
  assign s_1133 = 1'd1;
  assign s_1134 = s_1135[27];
  assign s_1135 = s_1136 - s_1143;
  assign s_1136 = s_1137;
  assign s_1137 = s_1138 | s_1142;
  assign s_1138 = s_1139 << s_1141;
  dq #(28, 1) dq_s_1139 (clk, s_1139, s_1140);
  assign s_1140 = s_1121?s_1124:s_1122;
  assign s_1141 = 1'd1;
  assign s_1142 = 1'd0;
  dq #(27, 19) dq_s_1143 (clk, s_1143, s_513);
  assign s_1144 = 1'd1;
  assign s_1145 = s_59 | s_1146;
  assign s_1146 = 1'd1;
  assign s_1147 = s_1148[27];
  assign s_1148 = s_1149 - s_1156;
  assign s_1149 = s_1150;
  assign s_1150 = s_1151 | s_1155;
  assign s_1151 = s_1152 << s_1154;
  dq #(28, 1) dq_s_1152 (clk, s_1152, s_1153);
  assign s_1153 = s_1134?s_1137:s_1135;
  assign s_1154 = 1'd1;
  assign s_1155 = 1'd0;
  dq #(27, 20) dq_s_1156 (clk, s_1156, s_513);
  assign s_1157 = 1'd1;
  assign s_1158 = s_56 | s_1159;
  assign s_1159 = 1'd1;
  assign s_1160 = s_1161[27];
  assign s_1161 = s_1162 - s_1169;
  assign s_1162 = s_1163;
  assign s_1163 = s_1164 | s_1168;
  assign s_1164 = s_1165 << s_1167;
  dq #(28, 1) dq_s_1165 (clk, s_1165, s_1166);
  assign s_1166 = s_1147?s_1150:s_1148;
  assign s_1167 = 1'd1;
  assign s_1168 = 1'd0;
  dq #(27, 21) dq_s_1169 (clk, s_1169, s_513);
  assign s_1170 = 1'd1;
  assign s_1171 = s_53 | s_1172;
  assign s_1172 = 1'd1;
  assign s_1173 = s_1174[27];
  assign s_1174 = s_1175 - s_1182;
  assign s_1175 = s_1176;
  assign s_1176 = s_1177 | s_1181;
  assign s_1177 = s_1178 << s_1180;
  dq #(28, 1) dq_s_1178 (clk, s_1178, s_1179);
  assign s_1179 = s_1160?s_1163:s_1161;
  assign s_1180 = 1'd1;
  assign s_1181 = 1'd0;
  dq #(27, 22) dq_s_1182 (clk, s_1182, s_513);
  assign s_1183 = 1'd1;
  assign s_1184 = s_50 | s_1185;
  assign s_1185 = 1'd1;
  assign s_1186 = s_1187[27];
  assign s_1187 = s_1188 - s_1195;
  assign s_1188 = s_1189;
  assign s_1189 = s_1190 | s_1194;
  assign s_1190 = s_1191 << s_1193;
  dq #(28, 1) dq_s_1191 (clk, s_1191, s_1192);
  assign s_1192 = s_1173?s_1176:s_1174;
  assign s_1193 = 1'd1;
  assign s_1194 = 1'd0;
  dq #(27, 23) dq_s_1195 (clk, s_1195, s_513);
  assign s_1196 = 1'd1;
  assign s_1197 = s_47 | s_1198;
  assign s_1198 = 1'd1;
  assign s_1199 = s_1200[27];
  assign s_1200 = s_1201 - s_1208;
  assign s_1201 = s_1202;
  assign s_1202 = s_1203 | s_1207;
  assign s_1203 = s_1204 << s_1206;
  dq #(28, 1) dq_s_1204 (clk, s_1204, s_1205);
  assign s_1205 = s_1186?s_1189:s_1187;
  assign s_1206 = 1'd1;
  assign s_1207 = 1'd0;
  dq #(27, 24) dq_s_1208 (clk, s_1208, s_513);
  assign s_1209 = 1'd1;
  assign s_1210 = s_44 | s_1211;
  assign s_1211 = 1'd1;
  assign s_1212 = s_1213[27];
  assign s_1213 = s_1214 - s_1221;
  assign s_1214 = s_1215;
  assign s_1215 = s_1216 | s_1220;
  assign s_1216 = s_1217 << s_1219;
  dq #(28, 1) dq_s_1217 (clk, s_1217, s_1218);
  assign s_1218 = s_1199?s_1202:s_1200;
  assign s_1219 = 1'd1;
  assign s_1220 = 1'd0;
  dq #(27, 25) dq_s_1221 (clk, s_1221, s_513);
  assign s_1222 = 1'd1;
  assign s_1223 = s_41 | s_1224;
  assign s_1224 = 1'd1;
  assign s_1225 = s_1226[27];
  assign s_1226 = s_1227 - s_1234;
  assign s_1227 = s_1228;
  assign s_1228 = s_1229 | s_1233;
  assign s_1229 = s_1230 << s_1232;
  dq #(28, 1) dq_s_1230 (clk, s_1230, s_1231);
  assign s_1231 = s_1212?s_1215:s_1213;
  assign s_1232 = 1'd1;
  assign s_1233 = 1'd0;
  dq #(27, 26) dq_s_1234 (clk, s_1234, s_513);
  dq #(10, 24) dq_s_1235 (clk, s_1235, s_1236);
  dq #(10, 1) dq_s_1236 (clk, s_1236, s_1237);
  assign s_1237 = s_1250?s_1238:s_1239;
  assign s_1238 = 1'd0;
  dq #(10, 1) dq_s_1239 (clk, s_1239, s_1240);
  assign s_1240 = s_1241 - s_1242;
  assign s_1241 = -10'd126;
  dq #(10, 1) dq_s_1242 (clk, s_1242, s_1243);
  assign s_1243 = s_1244 - s_1247;
  dq #(10, 1) dq_s_1244 (clk, s_1244, s_1245);
  assign s_1245 = s_1246 - s_144;
  dq #(10, 2) dq_s_1246 (clk, s_1246, s_505);
  dq #(10, 1) dq_s_1247 (clk, s_1247, s_1248);
  assign s_1248 = s_1249 - s_528;
  dq #(10, 2) dq_s_1249 (clk, s_1249, s_889);
  assign s_1250 = s_1239[9];
  dq #(10, 1) dq_s_1251 (clk, s_1251, s_1252);
  assign s_1252 = s_1610?s_1253:s_1604;
  dq #(6, 1) dq_s_1253 (clk, s_1253, s_1254);
  assign s_1254 = {s_1255,s_1598};
  assign s_1255 = s_1256 & s_1432;
  assign s_1256 = s_1257[4];
  assign s_1257 = {s_1258,s_1426};
  assign s_1258 = s_1259 & s_1348;
  assign s_1259 = s_1260[3];
  assign s_1260 = {s_1261,s_1342};
  assign s_1261 = s_1262 & s_1308;
  assign s_1262 = s_1263[2];
  assign s_1263 = {s_1264,s_1302};
  assign s_1264 = s_1265 & s_1290;
  assign s_1265 = s_1266[1];
  assign s_1266 = {s_1267,s_1286};
  assign s_1267 = s_1268 & s_1284;
  assign s_1268 = ~s_1269;
  assign s_1269 = s_1270[1];
  assign s_1270 = s_1271[3:2];
  assign s_1271 = s_1272[7:4];
  assign s_1272 = s_1273[15:8];
  assign s_1273 = s_1274[31:16];
  assign s_1274 = {s_1275,s_1283};
  assign s_1275 = {s_1276,s_1282};
  assign s_1276 = {s_1277,s_1281};
  assign s_1277 = {s_1278,s_1280};
  assign s_1278 = {s_37,s_1279};
  assign s_1279 = 1'd1;
  assign s_1280 = 1'd1;
  assign s_1281 = 1'd1;
  assign s_1282 = 1'd1;
  assign s_1283 = 1'd1;
  assign s_1284 = ~s_1285;
  assign s_1285 = s_1270[0];
  assign s_1286 = s_1287 & s_1289;
  assign s_1287 = ~s_1288;
  assign s_1288 = s_1270[1];
  assign s_1289 = s_1270[0];
  assign s_1290 = s_1291[1];
  assign s_1291 = {s_1292,s_1298};
  assign s_1292 = s_1293 & s_1296;
  assign s_1293 = ~s_1294;
  assign s_1294 = s_1295[1];
  assign s_1295 = s_1271[1:0];
  assign s_1296 = ~s_1297;
  assign s_1297 = s_1295[0];
  assign s_1298 = s_1299 & s_1301;
  assign s_1299 = ~s_1300;
  assign s_1300 = s_1295[1];
  assign s_1301 = s_1295[0];
  assign s_1302 = {s_1303,s_1305};
  assign s_1303 = s_1265 & s_1304;
  assign s_1304 = ~s_1290;
  assign s_1305 = s_1265?s_1306:s_1307;
  assign s_1306 = s_1291[0:0];
  assign s_1307 = s_1266[0:0];
  assign s_1308 = s_1309[2];
  assign s_1309 = {s_1310,s_1336};
  assign s_1310 = s_1311 & s_1324;
  assign s_1311 = s_1312[1];
  assign s_1312 = {s_1313,s_1320};
  assign s_1313 = s_1314 & s_1318;
  assign s_1314 = ~s_1315;
  assign s_1315 = s_1316[1];
  assign s_1316 = s_1317[3:2];
  assign s_1317 = s_1272[3:0];
  assign s_1318 = ~s_1319;
  assign s_1319 = s_1316[0];
  assign s_1320 = s_1321 & s_1323;
  assign s_1321 = ~s_1322;
  assign s_1322 = s_1316[1];
  assign s_1323 = s_1316[0];
  assign s_1324 = s_1325[1];
  assign s_1325 = {s_1326,s_1332};
  assign s_1326 = s_1327 & s_1330;
  assign s_1327 = ~s_1328;
  assign s_1328 = s_1329[1];
  assign s_1329 = s_1317[1:0];
  assign s_1330 = ~s_1331;
  assign s_1331 = s_1329[0];
  assign s_1332 = s_1333 & s_1335;
  assign s_1333 = ~s_1334;
  assign s_1334 = s_1329[1];
  assign s_1335 = s_1329[0];
  assign s_1336 = {s_1337,s_1339};
  assign s_1337 = s_1311 & s_1338;
  assign s_1338 = ~s_1324;
  assign s_1339 = s_1311?s_1340:s_1341;
  assign s_1340 = s_1325[0:0];
  assign s_1341 = s_1312[0:0];
  assign s_1342 = {s_1343,s_1345};
  assign s_1343 = s_1262 & s_1344;
  assign s_1344 = ~s_1308;
  assign s_1345 = s_1262?s_1346:s_1347;
  assign s_1346 = s_1309[1:0];
  assign s_1347 = s_1263[1:0];
  assign s_1348 = s_1349[3];
  assign s_1349 = {s_1350,s_1420};
  assign s_1350 = s_1351 & s_1386;
  assign s_1351 = s_1352[2];
  assign s_1352 = {s_1353,s_1380};
  assign s_1353 = s_1354 & s_1368;
  assign s_1354 = s_1355[1];
  assign s_1355 = {s_1356,s_1364};
  assign s_1356 = s_1357 & s_1362;
  assign s_1357 = ~s_1358;
  assign s_1358 = s_1359[1];
  assign s_1359 = s_1360[3:2];
  assign s_1360 = s_1361[7:4];
  assign s_1361 = s_1273[7:0];
  assign s_1362 = ~s_1363;
  assign s_1363 = s_1359[0];
  assign s_1364 = s_1365 & s_1367;
  assign s_1365 = ~s_1366;
  assign s_1366 = s_1359[1];
  assign s_1367 = s_1359[0];
  assign s_1368 = s_1369[1];
  assign s_1369 = {s_1370,s_1376};
  assign s_1370 = s_1371 & s_1374;
  assign s_1371 = ~s_1372;
  assign s_1372 = s_1373[1];
  assign s_1373 = s_1360[1:0];
  assign s_1374 = ~s_1375;
  assign s_1375 = s_1373[0];
  assign s_1376 = s_1377 & s_1379;
  assign s_1377 = ~s_1378;
  assign s_1378 = s_1373[1];
  assign s_1379 = s_1373[0];
  assign s_1380 = {s_1381,s_1383};
  assign s_1381 = s_1354 & s_1382;
  assign s_1382 = ~s_1368;
  assign s_1383 = s_1354?s_1384:s_1385;
  assign s_1384 = s_1369[0:0];
  assign s_1385 = s_1355[0:0];
  assign s_1386 = s_1387[2];
  assign s_1387 = {s_1388,s_1414};
  assign s_1388 = s_1389 & s_1402;
  assign s_1389 = s_1390[1];
  assign s_1390 = {s_1391,s_1398};
  assign s_1391 = s_1392 & s_1396;
  assign s_1392 = ~s_1393;
  assign s_1393 = s_1394[1];
  assign s_1394 = s_1395[3:2];
  assign s_1395 = s_1361[3:0];
  assign s_1396 = ~s_1397;
  assign s_1397 = s_1394[0];
  assign s_1398 = s_1399 & s_1401;
  assign s_1399 = ~s_1400;
  assign s_1400 = s_1394[1];
  assign s_1401 = s_1394[0];
  assign s_1402 = s_1403[1];
  assign s_1403 = {s_1404,s_1410};
  assign s_1404 = s_1405 & s_1408;
  assign s_1405 = ~s_1406;
  assign s_1406 = s_1407[1];
  assign s_1407 = s_1395[1:0];
  assign s_1408 = ~s_1409;
  assign s_1409 = s_1407[0];
  assign s_1410 = s_1411 & s_1413;
  assign s_1411 = ~s_1412;
  assign s_1412 = s_1407[1];
  assign s_1413 = s_1407[0];
  assign s_1414 = {s_1415,s_1417};
  assign s_1415 = s_1389 & s_1416;
  assign s_1416 = ~s_1402;
  assign s_1417 = s_1389?s_1418:s_1419;
  assign s_1418 = s_1403[0:0];
  assign s_1419 = s_1390[0:0];
  assign s_1420 = {s_1421,s_1423};
  assign s_1421 = s_1351 & s_1422;
  assign s_1422 = ~s_1386;
  assign s_1423 = s_1351?s_1424:s_1425;
  assign s_1424 = s_1387[1:0];
  assign s_1425 = s_1352[1:0];
  assign s_1426 = {s_1427,s_1429};
  assign s_1427 = s_1259 & s_1428;
  assign s_1428 = ~s_1348;
  assign s_1429 = s_1259?s_1430:s_1431;
  assign s_1430 = s_1349[2:0];
  assign s_1431 = s_1260[2:0];
  assign s_1432 = s_1433[4];
  assign s_1433 = {s_1434,s_1592};
  assign s_1434 = s_1435 & s_1514;
  assign s_1435 = s_1436[3];
  assign s_1436 = {s_1437,s_1508};
  assign s_1437 = s_1438 & s_1474;
  assign s_1438 = s_1439[2];
  assign s_1439 = {s_1440,s_1468};
  assign s_1440 = s_1441 & s_1456;
  assign s_1441 = s_1442[1];
  assign s_1442 = {s_1443,s_1452};
  assign s_1443 = s_1444 & s_1450;
  assign s_1444 = ~s_1445;
  assign s_1445 = s_1446[1];
  assign s_1446 = s_1447[3:2];
  assign s_1447 = s_1448[7:4];
  assign s_1448 = s_1449[15:8];
  assign s_1449 = s_1274[15:0];
  assign s_1450 = ~s_1451;
  assign s_1451 = s_1446[0];
  assign s_1452 = s_1453 & s_1455;
  assign s_1453 = ~s_1454;
  assign s_1454 = s_1446[1];
  assign s_1455 = s_1446[0];
  assign s_1456 = s_1457[1];
  assign s_1457 = {s_1458,s_1464};
  assign s_1458 = s_1459 & s_1462;
  assign s_1459 = ~s_1460;
  assign s_1460 = s_1461[1];
  assign s_1461 = s_1447[1:0];
  assign s_1462 = ~s_1463;
  assign s_1463 = s_1461[0];
  assign s_1464 = s_1465 & s_1467;
  assign s_1465 = ~s_1466;
  assign s_1466 = s_1461[1];
  assign s_1467 = s_1461[0];
  assign s_1468 = {s_1469,s_1471};
  assign s_1469 = s_1441 & s_1470;
  assign s_1470 = ~s_1456;
  assign s_1471 = s_1441?s_1472:s_1473;
  assign s_1472 = s_1457[0:0];
  assign s_1473 = s_1442[0:0];
  assign s_1474 = s_1475[2];
  assign s_1475 = {s_1476,s_1502};
  assign s_1476 = s_1477 & s_1490;
  assign s_1477 = s_1478[1];
  assign s_1478 = {s_1479,s_1486};
  assign s_1479 = s_1480 & s_1484;
  assign s_1480 = ~s_1481;
  assign s_1481 = s_1482[1];
  assign s_1482 = s_1483[3:2];
  assign s_1483 = s_1448[3:0];
  assign s_1484 = ~s_1485;
  assign s_1485 = s_1482[0];
  assign s_1486 = s_1487 & s_1489;
  assign s_1487 = ~s_1488;
  assign s_1488 = s_1482[1];
  assign s_1489 = s_1482[0];
  assign s_1490 = s_1491[1];
  assign s_1491 = {s_1492,s_1498};
  assign s_1492 = s_1493 & s_1496;
  assign s_1493 = ~s_1494;
  assign s_1494 = s_1495[1];
  assign s_1495 = s_1483[1:0];
  assign s_1496 = ~s_1497;
  assign s_1497 = s_1495[0];
  assign s_1498 = s_1499 & s_1501;
  assign s_1499 = ~s_1500;
  assign s_1500 = s_1495[1];
  assign s_1501 = s_1495[0];
  assign s_1502 = {s_1503,s_1505};
  assign s_1503 = s_1477 & s_1504;
  assign s_1504 = ~s_1490;
  assign s_1505 = s_1477?s_1506:s_1507;
  assign s_1506 = s_1491[0:0];
  assign s_1507 = s_1478[0:0];
  assign s_1508 = {s_1509,s_1511};
  assign s_1509 = s_1438 & s_1510;
  assign s_1510 = ~s_1474;
  assign s_1511 = s_1438?s_1512:s_1513;
  assign s_1512 = s_1475[1:0];
  assign s_1513 = s_1439[1:0];
  assign s_1514 = s_1515[3];
  assign s_1515 = {s_1516,s_1586};
  assign s_1516 = s_1517 & s_1552;
  assign s_1517 = s_1518[2];
  assign s_1518 = {s_1519,s_1546};
  assign s_1519 = s_1520 & s_1534;
  assign s_1520 = s_1521[1];
  assign s_1521 = {s_1522,s_1530};
  assign s_1522 = s_1523 & s_1528;
  assign s_1523 = ~s_1524;
  assign s_1524 = s_1525[1];
  assign s_1525 = s_1526[3:2];
  assign s_1526 = s_1527[7:4];
  assign s_1527 = s_1449[7:0];
  assign s_1528 = ~s_1529;
  assign s_1529 = s_1525[0];
  assign s_1530 = s_1531 & s_1533;
  assign s_1531 = ~s_1532;
  assign s_1532 = s_1525[1];
  assign s_1533 = s_1525[0];
  assign s_1534 = s_1535[1];
  assign s_1535 = {s_1536,s_1542};
  assign s_1536 = s_1537 & s_1540;
  assign s_1537 = ~s_1538;
  assign s_1538 = s_1539[1];
  assign s_1539 = s_1526[1:0];
  assign s_1540 = ~s_1541;
  assign s_1541 = s_1539[0];
  assign s_1542 = s_1543 & s_1545;
  assign s_1543 = ~s_1544;
  assign s_1544 = s_1539[1];
  assign s_1545 = s_1539[0];
  assign s_1546 = {s_1547,s_1549};
  assign s_1547 = s_1520 & s_1548;
  assign s_1548 = ~s_1534;
  assign s_1549 = s_1520?s_1550:s_1551;
  assign s_1550 = s_1535[0:0];
  assign s_1551 = s_1521[0:0];
  assign s_1552 = s_1553[2];
  assign s_1553 = {s_1554,s_1580};
  assign s_1554 = s_1555 & s_1568;
  assign s_1555 = s_1556[1];
  assign s_1556 = {s_1557,s_1564};
  assign s_1557 = s_1558 & s_1562;
  assign s_1558 = ~s_1559;
  assign s_1559 = s_1560[1];
  assign s_1560 = s_1561[3:2];
  assign s_1561 = s_1527[3:0];
  assign s_1562 = ~s_1563;
  assign s_1563 = s_1560[0];
  assign s_1564 = s_1565 & s_1567;
  assign s_1565 = ~s_1566;
  assign s_1566 = s_1560[1];
  assign s_1567 = s_1560[0];
  assign s_1568 = s_1569[1];
  assign s_1569 = {s_1570,s_1576};
  assign s_1570 = s_1571 & s_1574;
  assign s_1571 = ~s_1572;
  assign s_1572 = s_1573[1];
  assign s_1573 = s_1561[1:0];
  assign s_1574 = ~s_1575;
  assign s_1575 = s_1573[0];
  assign s_1576 = s_1577 & s_1579;
  assign s_1577 = ~s_1578;
  assign s_1578 = s_1573[1];
  assign s_1579 = s_1573[0];
  assign s_1580 = {s_1581,s_1583};
  assign s_1581 = s_1555 & s_1582;
  assign s_1582 = ~s_1568;
  assign s_1583 = s_1555?s_1584:s_1585;
  assign s_1584 = s_1569[0:0];
  assign s_1585 = s_1556[0:0];
  assign s_1586 = {s_1587,s_1589};
  assign s_1587 = s_1517 & s_1588;
  assign s_1588 = ~s_1552;
  assign s_1589 = s_1517?s_1590:s_1591;
  assign s_1590 = s_1553[1:0];
  assign s_1591 = s_1518[1:0];
  assign s_1592 = {s_1593,s_1595};
  assign s_1593 = s_1435 & s_1594;
  assign s_1594 = ~s_1514;
  assign s_1595 = s_1435?s_1596:s_1597;
  assign s_1596 = s_1515[2:0];
  assign s_1597 = s_1436[2:0];
  assign s_1598 = {s_1599,s_1601};
  assign s_1599 = s_1256 & s_1600;
  assign s_1600 = ~s_1432;
  assign s_1601 = s_1256?s_1602:s_1603;
  assign s_1602 = s_1433[3:0];
  assign s_1603 = s_1257[3:0];
  dq #(10, 25) dq_s_1604 (clk, s_1604, s_1605);
  assign s_1605 = s_1606 - s_1609;
  dq #(10, 1) dq_s_1606 (clk, s_1606, s_1607);
  assign s_1607 = s_1608 + s_1236;
  dq #(10, 2) dq_s_1608 (clk, s_1608, s_1242);
  assign s_1609 = -10'd126;
  assign s_1610 = s_1611 <= s_1612;
  assign s_1611 = s_1253;
  dq #(10, 25) dq_s_1612 (clk, s_1612, s_1605);
  assign s_1613 = 2'd3;
  assign s_1614 = 1'd1;
  dq #(24, 1) dq_s_1615 (clk, s_1615, s_32);
  assign s_1616 = s_1617 & s_1619;
  dq #(1, 1) dq_s_1617 (clk, s_1617, s_1618);
  assign s_1618 = s_34[2];
  assign s_1619 = s_1620 | s_1631;
  assign s_1620 = s_1621 | s_1623;
  dq #(1, 1) dq_s_1621 (clk, s_1621, s_1622);
  assign s_1622 = s_34[1];
  dq #(1, 1) dq_s_1623 (clk, s_1623, s_1624);
  assign s_1624 = s_1625 | s_1626;
  assign s_1625 = s_34[0];
  dq #(1, 4) dq_s_1626 (clk, s_1626, s_1627);
  assign s_1627 = s_1628 != s_1630;
  dq #(28, 1) dq_s_1628 (clk, s_1628, s_1629);
  assign s_1629 = s_1225?s_1228:s_1226;
  assign s_1630 = 1'd0;
  dq #(1, 1) dq_s_1631 (clk, s_1631, s_1632);
  assign s_1632 = s_32[0];
  assign s_1633 = s_28[23:0];
  assign s_1634 = s_28[24];
  dq #(1, 36) dq_s_1635 (clk, s_1635, s_1636);
  assign s_1636 = s_1637 & s_1639;
  assign s_1637 = s_523 == s_1638;
  assign s_1638 = 8'd128;
  assign s_1639 = s_527 == s_1640;
  assign s_1640 = 23'd0;
  assign s_1641 = {s_1642,s_1653};
  assign s_1642 = {s_1643,s_1644};
  dq #(1, 36) dq_s_1643 (clk, s_1643, s_3);
  assign s_1644 = s_1645 + s_1652;
  assign s_1645 = s_1646[7:0];
  dq #(10, 1) dq_s_1646 (clk, s_1646, s_1647);
  assign s_1647 = s_1648 + s_1634;
  dq #(10, 1) dq_s_1648 (clk, s_1648, s_1649);
  dq #(10, 1) dq_s_1649 (clk, s_1649, s_1650);
  assign s_1650 = s_1651 - s_1251;
  dq #(10, 26) dq_s_1651 (clk, s_1651, s_1606);
  assign s_1652 = 7'd127;
  assign s_1653 = s_23[22:0];
  assign s_1654 = s_1655 & s_1657;
  assign s_1655 = s_1645 == s_1656;
  assign s_1656 = -8'd126;
  assign s_1657 = ~s_1658;
  assign s_1658 = s_23[23];
  assign s_1659 = s_23 == s_1660;
  assign s_1660 = 24'd0;
  assign s_1661 = s_1677?s_1662:s_1663;
  assign s_1662 = 1'd0;
  assign s_1663 = s_1664 | s_1673;
  assign s_1664 = s_1665 | s_1667;
  assign s_1665 = $signed(s_1646) > $signed(s_1666);
  assign s_1666 = 9'd127;
  dq #(1, 36) dq_s_1667 (clk, s_1667, s_1668);
  assign s_1668 = s_1669 & s_1671;
  assign s_1669 = s_139 == s_1670;
  assign s_1670 = 8'd128;
  assign s_1671 = s_143 == s_1672;
  assign s_1672 = 23'd0;
  dq #(1, 32) dq_s_1673 (clk, s_1673, s_1674);
  dq #(1, 1) dq_s_1674 (clk, s_1674, s_1675);
  assign s_1675 = s_513 == s_1676;
  assign s_1676 = 1'd0;
  dq #(1, 36) dq_s_1677 (clk, s_1677, s_1636);
  dq #(1, 36) dq_s_1678 (clk, s_1678, s_1679);
  assign s_1679 = s_1680 | s_1691;
  assign s_1680 = s_1681 | s_1686;
  assign s_1681 = s_1682 & s_1684;
  assign s_1682 = s_139 == s_1683;
  assign s_1683 = 8'd128;
  assign s_1684 = s_143 != s_1685;
  assign s_1685 = 23'd0;
  assign s_1686 = s_1687 & s_1689;
  assign s_1687 = s_523 == s_1688;
  assign s_1688 = 8'd128;
  assign s_1689 = s_527 != s_1690;
  assign s_1690 = 23'd0;
  assign s_1691 = s_1668 & s_1636;
  assign div_z = s_0;
endmodule
