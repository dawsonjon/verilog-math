module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module unsigned_int_to_single(clk, unsigned_int_to_single_a, unsigned_int_to_single_z);
  input clk;
  input [31:0] unsigned_int_to_single_a;
  output [31:0] unsigned_int_to_single_z;
  wire [31:0] s_0;
  wire [31:0] s_1;
  wire [31:0] s_2;
  wire [0:0] s_3;
  wire [30:0] s_4;
  wire [31:0] s_5;
  wire [31:0] s_6;
  wire [31:0] s_7;
  wire [30:0] s_8;
  wire [31:0] s_9;
  wire [31:0] s_10;
  wire [31:0] s_11;
  wire [30:0] s_12;
  wire [31:0] s_13;
  wire [31:0] s_14;
  wire [8:0] s_15;
  wire [8:0] s_16;
  wire [7:0] s_17;
  wire [22:0] s_18;
  wire [23:0] s_19;
  wire [23:0] s_20;
  wire [23:0] s_21;
  wire [24:0] s_22;
  wire [24:0] s_23;
  wire [24:0] s_24;
  wire [24:0] s_25;
  wire [23:0] s_26;
  wire [31:0] s_27;
  wire [31:0] s_28;
  wire [31:0] s_29;
  wire [31:0] s_30;
  wire [31:0] s_31;
  wire [5:0] s_32;
  wire [5:0] s_33;
  wire [0:0] s_34;
  wire [0:0] s_35;
  wire [4:0] s_36;
  wire [0:0] s_37;
  wire [0:0] s_38;
  wire [3:0] s_39;
  wire [0:0] s_40;
  wire [0:0] s_41;
  wire [2:0] s_42;
  wire [0:0] s_43;
  wire [0:0] s_44;
  wire [1:0] s_45;
  wire [0:0] s_46;
  wire [0:0] s_47;
  wire [0:0] s_48;
  wire [1:0] s_49;
  wire [3:0] s_50;
  wire [7:0] s_51;
  wire [15:0] s_52;
  wire [0:0] s_53;
  wire [0:0] s_54;
  wire [0:0] s_55;
  wire [0:0] s_56;
  wire [0:0] s_57;
  wire [0:0] s_58;
  wire [0:0] s_59;
  wire [1:0] s_60;
  wire [0:0] s_61;
  wire [0:0] s_62;
  wire [0:0] s_63;
  wire [1:0] s_64;
  wire [0:0] s_65;
  wire [0:0] s_66;
  wire [0:0] s_67;
  wire [0:0] s_68;
  wire [0:0] s_69;
  wire [0:0] s_70;
  wire [1:0] s_71;
  wire [0:0] s_72;
  wire [0:0] s_73;
  wire [0:0] s_74;
  wire [0:0] s_75;
  wire [0:0] s_76;
  wire [0:0] s_77;
  wire [2:0] s_78;
  wire [0:0] s_79;
  wire [0:0] s_80;
  wire [1:0] s_81;
  wire [0:0] s_82;
  wire [0:0] s_83;
  wire [0:0] s_84;
  wire [1:0] s_85;
  wire [3:0] s_86;
  wire [0:0] s_87;
  wire [0:0] s_88;
  wire [0:0] s_89;
  wire [0:0] s_90;
  wire [0:0] s_91;
  wire [0:0] s_92;
  wire [0:0] s_93;
  wire [1:0] s_94;
  wire [0:0] s_95;
  wire [0:0] s_96;
  wire [0:0] s_97;
  wire [1:0] s_98;
  wire [0:0] s_99;
  wire [0:0] s_100;
  wire [0:0] s_101;
  wire [0:0] s_102;
  wire [0:0] s_103;
  wire [0:0] s_104;
  wire [1:0] s_105;
  wire [0:0] s_106;
  wire [0:0] s_107;
  wire [0:0] s_108;
  wire [0:0] s_109;
  wire [0:0] s_110;
  wire [2:0] s_111;
  wire [0:0] s_112;
  wire [0:0] s_113;
  wire [1:0] s_114;
  wire [1:0] s_115;
  wire [1:0] s_116;
  wire [0:0] s_117;
  wire [3:0] s_118;
  wire [0:0] s_119;
  wire [0:0] s_120;
  wire [2:0] s_121;
  wire [0:0] s_122;
  wire [0:0] s_123;
  wire [1:0] s_124;
  wire [0:0] s_125;
  wire [0:0] s_126;
  wire [0:0] s_127;
  wire [1:0] s_128;
  wire [3:0] s_129;
  wire [7:0] s_130;
  wire [0:0] s_131;
  wire [0:0] s_132;
  wire [0:0] s_133;
  wire [0:0] s_134;
  wire [0:0] s_135;
  wire [0:0] s_136;
  wire [0:0] s_137;
  wire [1:0] s_138;
  wire [0:0] s_139;
  wire [0:0] s_140;
  wire [0:0] s_141;
  wire [1:0] s_142;
  wire [0:0] s_143;
  wire [0:0] s_144;
  wire [0:0] s_145;
  wire [0:0] s_146;
  wire [0:0] s_147;
  wire [0:0] s_148;
  wire [1:0] s_149;
  wire [0:0] s_150;
  wire [0:0] s_151;
  wire [0:0] s_152;
  wire [0:0] s_153;
  wire [0:0] s_154;
  wire [0:0] s_155;
  wire [2:0] s_156;
  wire [0:0] s_157;
  wire [0:0] s_158;
  wire [1:0] s_159;
  wire [0:0] s_160;
  wire [0:0] s_161;
  wire [0:0] s_162;
  wire [1:0] s_163;
  wire [3:0] s_164;
  wire [0:0] s_165;
  wire [0:0] s_166;
  wire [0:0] s_167;
  wire [0:0] s_168;
  wire [0:0] s_169;
  wire [0:0] s_170;
  wire [0:0] s_171;
  wire [1:0] s_172;
  wire [0:0] s_173;
  wire [0:0] s_174;
  wire [0:0] s_175;
  wire [1:0] s_176;
  wire [0:0] s_177;
  wire [0:0] s_178;
  wire [0:0] s_179;
  wire [0:0] s_180;
  wire [0:0] s_181;
  wire [0:0] s_182;
  wire [1:0] s_183;
  wire [0:0] s_184;
  wire [0:0] s_185;
  wire [0:0] s_186;
  wire [0:0] s_187;
  wire [0:0] s_188;
  wire [2:0] s_189;
  wire [0:0] s_190;
  wire [0:0] s_191;
  wire [1:0] s_192;
  wire [1:0] s_193;
  wire [1:0] s_194;
  wire [3:0] s_195;
  wire [0:0] s_196;
  wire [0:0] s_197;
  wire [2:0] s_198;
  wire [2:0] s_199;
  wire [2:0] s_200;
  wire [0:0] s_201;
  wire [4:0] s_202;
  wire [0:0] s_203;
  wire [0:0] s_204;
  wire [3:0] s_205;
  wire [0:0] s_206;
  wire [0:0] s_207;
  wire [2:0] s_208;
  wire [0:0] s_209;
  wire [0:0] s_210;
  wire [1:0] s_211;
  wire [0:0] s_212;
  wire [0:0] s_213;
  wire [0:0] s_214;
  wire [1:0] s_215;
  wire [3:0] s_216;
  wire [7:0] s_217;
  wire [15:0] s_218;
  wire [0:0] s_219;
  wire [0:0] s_220;
  wire [0:0] s_221;
  wire [0:0] s_222;
  wire [0:0] s_223;
  wire [0:0] s_224;
  wire [0:0] s_225;
  wire [1:0] s_226;
  wire [0:0] s_227;
  wire [0:0] s_228;
  wire [0:0] s_229;
  wire [1:0] s_230;
  wire [0:0] s_231;
  wire [0:0] s_232;
  wire [0:0] s_233;
  wire [0:0] s_234;
  wire [0:0] s_235;
  wire [0:0] s_236;
  wire [1:0] s_237;
  wire [0:0] s_238;
  wire [0:0] s_239;
  wire [0:0] s_240;
  wire [0:0] s_241;
  wire [0:0] s_242;
  wire [0:0] s_243;
  wire [2:0] s_244;
  wire [0:0] s_245;
  wire [0:0] s_246;
  wire [1:0] s_247;
  wire [0:0] s_248;
  wire [0:0] s_249;
  wire [0:0] s_250;
  wire [1:0] s_251;
  wire [3:0] s_252;
  wire [0:0] s_253;
  wire [0:0] s_254;
  wire [0:0] s_255;
  wire [0:0] s_256;
  wire [0:0] s_257;
  wire [0:0] s_258;
  wire [0:0] s_259;
  wire [1:0] s_260;
  wire [0:0] s_261;
  wire [0:0] s_262;
  wire [0:0] s_263;
  wire [1:0] s_264;
  wire [0:0] s_265;
  wire [0:0] s_266;
  wire [0:0] s_267;
  wire [0:0] s_268;
  wire [0:0] s_269;
  wire [0:0] s_270;
  wire [1:0] s_271;
  wire [0:0] s_272;
  wire [0:0] s_273;
  wire [0:0] s_274;
  wire [0:0] s_275;
  wire [0:0] s_276;
  wire [2:0] s_277;
  wire [0:0] s_278;
  wire [0:0] s_279;
  wire [1:0] s_280;
  wire [1:0] s_281;
  wire [1:0] s_282;
  wire [0:0] s_283;
  wire [3:0] s_284;
  wire [0:0] s_285;
  wire [0:0] s_286;
  wire [2:0] s_287;
  wire [0:0] s_288;
  wire [0:0] s_289;
  wire [1:0] s_290;
  wire [0:0] s_291;
  wire [0:0] s_292;
  wire [0:0] s_293;
  wire [1:0] s_294;
  wire [3:0] s_295;
  wire [7:0] s_296;
  wire [0:0] s_297;
  wire [0:0] s_298;
  wire [0:0] s_299;
  wire [0:0] s_300;
  wire [0:0] s_301;
  wire [0:0] s_302;
  wire [0:0] s_303;
  wire [1:0] s_304;
  wire [0:0] s_305;
  wire [0:0] s_306;
  wire [0:0] s_307;
  wire [1:0] s_308;
  wire [0:0] s_309;
  wire [0:0] s_310;
  wire [0:0] s_311;
  wire [0:0] s_312;
  wire [0:0] s_313;
  wire [0:0] s_314;
  wire [1:0] s_315;
  wire [0:0] s_316;
  wire [0:0] s_317;
  wire [0:0] s_318;
  wire [0:0] s_319;
  wire [0:0] s_320;
  wire [0:0] s_321;
  wire [2:0] s_322;
  wire [0:0] s_323;
  wire [0:0] s_324;
  wire [1:0] s_325;
  wire [0:0] s_326;
  wire [0:0] s_327;
  wire [0:0] s_328;
  wire [1:0] s_329;
  wire [3:0] s_330;
  wire [0:0] s_331;
  wire [0:0] s_332;
  wire [0:0] s_333;
  wire [0:0] s_334;
  wire [0:0] s_335;
  wire [0:0] s_336;
  wire [0:0] s_337;
  wire [1:0] s_338;
  wire [0:0] s_339;
  wire [0:0] s_340;
  wire [0:0] s_341;
  wire [1:0] s_342;
  wire [0:0] s_343;
  wire [0:0] s_344;
  wire [0:0] s_345;
  wire [0:0] s_346;
  wire [0:0] s_347;
  wire [0:0] s_348;
  wire [1:0] s_349;
  wire [0:0] s_350;
  wire [0:0] s_351;
  wire [0:0] s_352;
  wire [0:0] s_353;
  wire [0:0] s_354;
  wire [2:0] s_355;
  wire [0:0] s_356;
  wire [0:0] s_357;
  wire [1:0] s_358;
  wire [1:0] s_359;
  wire [1:0] s_360;
  wire [3:0] s_361;
  wire [0:0] s_362;
  wire [0:0] s_363;
  wire [2:0] s_364;
  wire [2:0] s_365;
  wire [2:0] s_366;
  wire [4:0] s_367;
  wire [0:0] s_368;
  wire [0:0] s_369;
  wire [3:0] s_370;
  wire [3:0] s_371;
  wire [3:0] s_372;
  wire [0:0] s_373;
  wire [23:0] s_374;
  wire [0:0] s_375;
  wire [0:0] s_376;
  wire [0:0] s_377;
  wire [0:0] s_378;
  wire [0:0] s_379;
  wire [0:0] s_380;
  wire [0:0] s_381;
  wire [0:0] s_382;
  wire [0:0] s_383;
  wire [5:0] s_384;
  wire [0:0] s_385;
  wire [0:0] s_386;
  wire [0:0] s_387;
  wire [23:0] s_388;
  wire [0:0] s_389;
  wire [31:0] s_390;
  wire [8:0] s_391;
  wire [7:0] s_392;
  wire [7:0] s_393;
  wire [7:0] s_394;
  wire [7:0] s_395;
  wire [7:0] s_396;
  wire [7:0] s_397;
  wire [6:0] s_398;
  wire [22:0] s_399;
  wire [0:0] s_400;
  wire [0:0] s_401;
  wire [7:0] s_402;
  wire [0:0] s_403;
  wire [0:0] s_404;
  wire [0:0] s_405;
  wire [23:0] s_406;
  wire [0:0] s_407;
  wire [0:0] s_408;

  assign s_0 = s_408?s_1:s_5;
  dq #(32, 5) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_4};
  assign s_3 = 1'd0;
  assign s_4 = 31'd2143289344;
  assign s_5 = s_407?s_6:s_9;
  dq #(32, 5) dq_s_6 (clk, s_6, s_7);
  assign s_7 = {s_3,s_8};
  assign s_8 = 31'd2139095040;
  assign s_9 = s_405?s_10:s_13;
  dq #(32, 5) dq_s_10 (clk, s_10, s_11);
  assign s_11 = {s_3,s_12};
  assign s_12 = 31'd0;
  assign s_13 = s_400?s_14:s_390;
  assign s_14 = {s_15,s_18};
  dq #(9, 5) dq_s_15 (clk, s_15, s_16);
  assign s_16 = {s_3,s_17};
  assign s_17 = 8'd0;
  assign s_18 = s_19[22:0];
  dq #(24, 1) dq_s_19 (clk, s_19, s_20);
  assign s_20 = s_389?s_21:s_388;
  assign s_21 = s_22[24:1];
  assign s_22 = s_375?s_23:s_374;
  dq #(25, 1) dq_s_23 (clk, s_23, s_24);
  assign s_24 = s_25 + s_373;
  assign s_25 = s_26;
  assign s_26 = s_27[31:8];
  dq #(32, 1) dq_s_27 (clk, s_27, s_28);
  assign s_28 = s_29 << s_32;
  dq #(32, 1) dq_s_29 (clk, s_29, s_30);
  dq #(32, 1) dq_s_30 (clk, s_30, s_31);
  assign s_31 = unsigned_int_to_single_a;
  dq #(6, 1) dq_s_32 (clk, s_32, s_33);
  assign s_33 = {s_34,s_367};
  assign s_34 = s_35 & s_201;
  assign s_35 = s_36[4];
  assign s_36 = {s_37,s_195};
  assign s_37 = s_38 & s_117;
  assign s_38 = s_39[3];
  assign s_39 = {s_40,s_111};
  assign s_40 = s_41 & s_77;
  assign s_41 = s_42[2];
  assign s_42 = {s_43,s_71};
  assign s_43 = s_44 & s_59;
  assign s_44 = s_45[1];
  assign s_45 = {s_46,s_55};
  assign s_46 = s_47 & s_53;
  assign s_47 = ~s_48;
  assign s_48 = s_49[1];
  assign s_49 = s_50[3:2];
  assign s_50 = s_51[7:4];
  assign s_51 = s_52[15:8];
  assign s_52 = s_30[31:16];
  assign s_53 = ~s_54;
  assign s_54 = s_49[0];
  assign s_55 = s_56 & s_58;
  assign s_56 = ~s_57;
  assign s_57 = s_49[1];
  assign s_58 = s_49[0];
  assign s_59 = s_60[1];
  assign s_60 = {s_61,s_67};
  assign s_61 = s_62 & s_65;
  assign s_62 = ~s_63;
  assign s_63 = s_64[1];
  assign s_64 = s_50[1:0];
  assign s_65 = ~s_66;
  assign s_66 = s_64[0];
  assign s_67 = s_68 & s_70;
  assign s_68 = ~s_69;
  assign s_69 = s_64[1];
  assign s_70 = s_64[0];
  assign s_71 = {s_72,s_74};
  assign s_72 = s_44 & s_73;
  assign s_73 = ~s_59;
  assign s_74 = s_44?s_75:s_76;
  assign s_75 = s_60[0:0];
  assign s_76 = s_45[0:0];
  assign s_77 = s_78[2];
  assign s_78 = {s_79,s_105};
  assign s_79 = s_80 & s_93;
  assign s_80 = s_81[1];
  assign s_81 = {s_82,s_89};
  assign s_82 = s_83 & s_87;
  assign s_83 = ~s_84;
  assign s_84 = s_85[1];
  assign s_85 = s_86[3:2];
  assign s_86 = s_51[3:0];
  assign s_87 = ~s_88;
  assign s_88 = s_85[0];
  assign s_89 = s_90 & s_92;
  assign s_90 = ~s_91;
  assign s_91 = s_85[1];
  assign s_92 = s_85[0];
  assign s_93 = s_94[1];
  assign s_94 = {s_95,s_101};
  assign s_95 = s_96 & s_99;
  assign s_96 = ~s_97;
  assign s_97 = s_98[1];
  assign s_98 = s_86[1:0];
  assign s_99 = ~s_100;
  assign s_100 = s_98[0];
  assign s_101 = s_102 & s_104;
  assign s_102 = ~s_103;
  assign s_103 = s_98[1];
  assign s_104 = s_98[0];
  assign s_105 = {s_106,s_108};
  assign s_106 = s_80 & s_107;
  assign s_107 = ~s_93;
  assign s_108 = s_80?s_109:s_110;
  assign s_109 = s_94[0:0];
  assign s_110 = s_81[0:0];
  assign s_111 = {s_112,s_114};
  assign s_112 = s_41 & s_113;
  assign s_113 = ~s_77;
  assign s_114 = s_41?s_115:s_116;
  assign s_115 = s_78[1:0];
  assign s_116 = s_42[1:0];
  assign s_117 = s_118[3];
  assign s_118 = {s_119,s_189};
  assign s_119 = s_120 & s_155;
  assign s_120 = s_121[2];
  assign s_121 = {s_122,s_149};
  assign s_122 = s_123 & s_137;
  assign s_123 = s_124[1];
  assign s_124 = {s_125,s_133};
  assign s_125 = s_126 & s_131;
  assign s_126 = ~s_127;
  assign s_127 = s_128[1];
  assign s_128 = s_129[3:2];
  assign s_129 = s_130[7:4];
  assign s_130 = s_52[7:0];
  assign s_131 = ~s_132;
  assign s_132 = s_128[0];
  assign s_133 = s_134 & s_136;
  assign s_134 = ~s_135;
  assign s_135 = s_128[1];
  assign s_136 = s_128[0];
  assign s_137 = s_138[1];
  assign s_138 = {s_139,s_145};
  assign s_139 = s_140 & s_143;
  assign s_140 = ~s_141;
  assign s_141 = s_142[1];
  assign s_142 = s_129[1:0];
  assign s_143 = ~s_144;
  assign s_144 = s_142[0];
  assign s_145 = s_146 & s_148;
  assign s_146 = ~s_147;
  assign s_147 = s_142[1];
  assign s_148 = s_142[0];
  assign s_149 = {s_150,s_152};
  assign s_150 = s_123 & s_151;
  assign s_151 = ~s_137;
  assign s_152 = s_123?s_153:s_154;
  assign s_153 = s_138[0:0];
  assign s_154 = s_124[0:0];
  assign s_155 = s_156[2];
  assign s_156 = {s_157,s_183};
  assign s_157 = s_158 & s_171;
  assign s_158 = s_159[1];
  assign s_159 = {s_160,s_167};
  assign s_160 = s_161 & s_165;
  assign s_161 = ~s_162;
  assign s_162 = s_163[1];
  assign s_163 = s_164[3:2];
  assign s_164 = s_130[3:0];
  assign s_165 = ~s_166;
  assign s_166 = s_163[0];
  assign s_167 = s_168 & s_170;
  assign s_168 = ~s_169;
  assign s_169 = s_163[1];
  assign s_170 = s_163[0];
  assign s_171 = s_172[1];
  assign s_172 = {s_173,s_179};
  assign s_173 = s_174 & s_177;
  assign s_174 = ~s_175;
  assign s_175 = s_176[1];
  assign s_176 = s_164[1:0];
  assign s_177 = ~s_178;
  assign s_178 = s_176[0];
  assign s_179 = s_180 & s_182;
  assign s_180 = ~s_181;
  assign s_181 = s_176[1];
  assign s_182 = s_176[0];
  assign s_183 = {s_184,s_186};
  assign s_184 = s_158 & s_185;
  assign s_185 = ~s_171;
  assign s_186 = s_158?s_187:s_188;
  assign s_187 = s_172[0:0];
  assign s_188 = s_159[0:0];
  assign s_189 = {s_190,s_192};
  assign s_190 = s_120 & s_191;
  assign s_191 = ~s_155;
  assign s_192 = s_120?s_193:s_194;
  assign s_193 = s_156[1:0];
  assign s_194 = s_121[1:0];
  assign s_195 = {s_196,s_198};
  assign s_196 = s_38 & s_197;
  assign s_197 = ~s_117;
  assign s_198 = s_38?s_199:s_200;
  assign s_199 = s_118[2:0];
  assign s_200 = s_39[2:0];
  assign s_201 = s_202[4];
  assign s_202 = {s_203,s_361};
  assign s_203 = s_204 & s_283;
  assign s_204 = s_205[3];
  assign s_205 = {s_206,s_277};
  assign s_206 = s_207 & s_243;
  assign s_207 = s_208[2];
  assign s_208 = {s_209,s_237};
  assign s_209 = s_210 & s_225;
  assign s_210 = s_211[1];
  assign s_211 = {s_212,s_221};
  assign s_212 = s_213 & s_219;
  assign s_213 = ~s_214;
  assign s_214 = s_215[1];
  assign s_215 = s_216[3:2];
  assign s_216 = s_217[7:4];
  assign s_217 = s_218[15:8];
  assign s_218 = s_30[15:0];
  assign s_219 = ~s_220;
  assign s_220 = s_215[0];
  assign s_221 = s_222 & s_224;
  assign s_222 = ~s_223;
  assign s_223 = s_215[1];
  assign s_224 = s_215[0];
  assign s_225 = s_226[1];
  assign s_226 = {s_227,s_233};
  assign s_227 = s_228 & s_231;
  assign s_228 = ~s_229;
  assign s_229 = s_230[1];
  assign s_230 = s_216[1:0];
  assign s_231 = ~s_232;
  assign s_232 = s_230[0];
  assign s_233 = s_234 & s_236;
  assign s_234 = ~s_235;
  assign s_235 = s_230[1];
  assign s_236 = s_230[0];
  assign s_237 = {s_238,s_240};
  assign s_238 = s_210 & s_239;
  assign s_239 = ~s_225;
  assign s_240 = s_210?s_241:s_242;
  assign s_241 = s_226[0:0];
  assign s_242 = s_211[0:0];
  assign s_243 = s_244[2];
  assign s_244 = {s_245,s_271};
  assign s_245 = s_246 & s_259;
  assign s_246 = s_247[1];
  assign s_247 = {s_248,s_255};
  assign s_248 = s_249 & s_253;
  assign s_249 = ~s_250;
  assign s_250 = s_251[1];
  assign s_251 = s_252[3:2];
  assign s_252 = s_217[3:0];
  assign s_253 = ~s_254;
  assign s_254 = s_251[0];
  assign s_255 = s_256 & s_258;
  assign s_256 = ~s_257;
  assign s_257 = s_251[1];
  assign s_258 = s_251[0];
  assign s_259 = s_260[1];
  assign s_260 = {s_261,s_267};
  assign s_261 = s_262 & s_265;
  assign s_262 = ~s_263;
  assign s_263 = s_264[1];
  assign s_264 = s_252[1:0];
  assign s_265 = ~s_266;
  assign s_266 = s_264[0];
  assign s_267 = s_268 & s_270;
  assign s_268 = ~s_269;
  assign s_269 = s_264[1];
  assign s_270 = s_264[0];
  assign s_271 = {s_272,s_274};
  assign s_272 = s_246 & s_273;
  assign s_273 = ~s_259;
  assign s_274 = s_246?s_275:s_276;
  assign s_275 = s_260[0:0];
  assign s_276 = s_247[0:0];
  assign s_277 = {s_278,s_280};
  assign s_278 = s_207 & s_279;
  assign s_279 = ~s_243;
  assign s_280 = s_207?s_281:s_282;
  assign s_281 = s_244[1:0];
  assign s_282 = s_208[1:0];
  assign s_283 = s_284[3];
  assign s_284 = {s_285,s_355};
  assign s_285 = s_286 & s_321;
  assign s_286 = s_287[2];
  assign s_287 = {s_288,s_315};
  assign s_288 = s_289 & s_303;
  assign s_289 = s_290[1];
  assign s_290 = {s_291,s_299};
  assign s_291 = s_292 & s_297;
  assign s_292 = ~s_293;
  assign s_293 = s_294[1];
  assign s_294 = s_295[3:2];
  assign s_295 = s_296[7:4];
  assign s_296 = s_218[7:0];
  assign s_297 = ~s_298;
  assign s_298 = s_294[0];
  assign s_299 = s_300 & s_302;
  assign s_300 = ~s_301;
  assign s_301 = s_294[1];
  assign s_302 = s_294[0];
  assign s_303 = s_304[1];
  assign s_304 = {s_305,s_311};
  assign s_305 = s_306 & s_309;
  assign s_306 = ~s_307;
  assign s_307 = s_308[1];
  assign s_308 = s_295[1:0];
  assign s_309 = ~s_310;
  assign s_310 = s_308[0];
  assign s_311 = s_312 & s_314;
  assign s_312 = ~s_313;
  assign s_313 = s_308[1];
  assign s_314 = s_308[0];
  assign s_315 = {s_316,s_318};
  assign s_316 = s_289 & s_317;
  assign s_317 = ~s_303;
  assign s_318 = s_289?s_319:s_320;
  assign s_319 = s_304[0:0];
  assign s_320 = s_290[0:0];
  assign s_321 = s_322[2];
  assign s_322 = {s_323,s_349};
  assign s_323 = s_324 & s_337;
  assign s_324 = s_325[1];
  assign s_325 = {s_326,s_333};
  assign s_326 = s_327 & s_331;
  assign s_327 = ~s_328;
  assign s_328 = s_329[1];
  assign s_329 = s_330[3:2];
  assign s_330 = s_296[3:0];
  assign s_331 = ~s_332;
  assign s_332 = s_329[0];
  assign s_333 = s_334 & s_336;
  assign s_334 = ~s_335;
  assign s_335 = s_329[1];
  assign s_336 = s_329[0];
  assign s_337 = s_338[1];
  assign s_338 = {s_339,s_345};
  assign s_339 = s_340 & s_343;
  assign s_340 = ~s_341;
  assign s_341 = s_342[1];
  assign s_342 = s_330[1:0];
  assign s_343 = ~s_344;
  assign s_344 = s_342[0];
  assign s_345 = s_346 & s_348;
  assign s_346 = ~s_347;
  assign s_347 = s_342[1];
  assign s_348 = s_342[0];
  assign s_349 = {s_350,s_352};
  assign s_350 = s_324 & s_351;
  assign s_351 = ~s_337;
  assign s_352 = s_324?s_353:s_354;
  assign s_353 = s_338[0:0];
  assign s_354 = s_325[0:0];
  assign s_355 = {s_356,s_358};
  assign s_356 = s_286 & s_357;
  assign s_357 = ~s_321;
  assign s_358 = s_286?s_359:s_360;
  assign s_359 = s_322[1:0];
  assign s_360 = s_287[1:0];
  assign s_361 = {s_362,s_364};
  assign s_362 = s_204 & s_363;
  assign s_363 = ~s_283;
  assign s_364 = s_204?s_365:s_366;
  assign s_365 = s_284[2:0];
  assign s_366 = s_205[2:0];
  assign s_367 = {s_368,s_370};
  assign s_368 = s_35 & s_369;
  assign s_369 = ~s_201;
  assign s_370 = s_35?s_371:s_372;
  assign s_371 = s_202[3:0];
  assign s_372 = s_36[3:0];
  assign s_373 = 1'd1;
  dq #(24, 1) dq_s_374 (clk, s_374, s_26);
  assign s_375 = s_376 & s_378;
  dq #(1, 1) dq_s_376 (clk, s_376, s_377);
  assign s_377 = s_27[7];
  assign s_378 = s_379 | s_386;
  assign s_379 = s_380 | s_382;
  dq #(1, 1) dq_s_380 (clk, s_380, s_381);
  assign s_381 = s_27[6];
  dq #(1, 1) dq_s_382 (clk, s_382, s_383);
  assign s_383 = s_384 != s_385;
  assign s_384 = s_27[5:0];
  assign s_385 = 1'd0;
  dq #(1, 1) dq_s_386 (clk, s_386, s_387);
  assign s_387 = s_26[0];
  assign s_388 = s_22[23:0];
  assign s_389 = s_22[24];
  assign s_390 = {s_391,s_399};
  assign s_391 = {s_3,s_392};
  assign s_392 = s_393 + s_398;
  dq #(8, 1) dq_s_393 (clk, s_393, s_394);
  assign s_394 = s_395 + s_389;
  dq #(8, 2) dq_s_395 (clk, s_395, s_396);
  assign s_396 = s_397 - s_32;
  assign s_397 = 8'd31;
  assign s_398 = 7'd127;
  assign s_399 = s_19[22:0];
  assign s_400 = s_401 & s_403;
  assign s_401 = s_393 == s_402;
  assign s_402 = -8'd126;
  assign s_403 = ~s_404;
  assign s_404 = s_19[23];
  assign s_405 = s_19 == s_406;
  assign s_406 = 24'd0;
  assign s_407 = 1'd0;
  assign s_408 = 1'd0;
  assign unsigned_int_to_single_z = s_0;
endmodule
