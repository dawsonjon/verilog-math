module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module mul(clk, mul_a, mul_b, mul_z);
  input clk;
  input [31:0] mul_a;
  input [31:0] mul_b;
  output [31:0] mul_z;
  wire [31:0] s_0;
  wire [31:0] s_1;
  wire [31:0] s_2;
  wire [0:0] s_3;
  wire [0:0] s_4;
  wire [31:0] s_5;
  wire [0:0] s_6;
  wire [31:0] s_7;
  wire [30:0] s_8;
  wire [31:0] s_9;
  wire [31:0] s_10;
  wire [31:0] s_11;
  wire [30:0] s_12;
  wire [31:0] s_13;
  wire [31:0] s_14;
  wire [31:0] s_15;
  wire [30:0] s_16;
  wire [31:0] s_17;
  wire [31:0] s_18;
  wire [8:0] s_19;
  wire [8:0] s_20;
  wire [7:0] s_21;
  wire [22:0] s_22;
  wire [23:0] s_23;
  wire [23:0] s_24;
  wire [23:0] s_25;
  wire [24:0] s_26;
  wire [24:0] s_27;
  wire [24:0] s_28;
  wire [24:0] s_29;
  wire [23:0] s_30;
  wire [47:0] s_31;
  wire [47:0] s_32;
  wire [47:0] s_33;
  wire [47:0] s_34;
  wire [47:0] s_35;
  wire [47:0] s_36;
  wire [47:0] s_37;
  wire [23:0] s_38;
  wire [0:0] s_39;
  wire [0:0] s_40;
  wire [0:0] s_41;
  wire [0:0] s_42;
  wire [7:0] s_43;
  wire [7:0] s_44;
  wire [6:0] s_45;
  wire [7:0] s_46;
  wire [22:0] s_47;
  wire [47:0] s_48;
  wire [23:0] s_49;
  wire [0:0] s_50;
  wire [0:0] s_51;
  wire [0:0] s_52;
  wire [0:0] s_53;
  wire [7:0] s_54;
  wire [7:0] s_55;
  wire [6:0] s_56;
  wire [7:0] s_57;
  wire [22:0] s_58;
  wire [9:0] s_59;
  wire [0:0] s_60;
  wire [9:0] s_61;
  wire [9:0] s_62;
  wire [9:0] s_63;
  wire [9:0] s_64;
  wire [9:0] s_65;
  wire [7:0] s_66;
  wire [7:0] s_67;
  wire [9:0] s_68;
  wire [7:0] s_69;
  wire [7:0] s_70;
  wire [0:0] s_71;
  wire [0:0] s_72;
  wire [9:0] s_73;
  wire [9:0] s_74;
  wire [6:0] s_75;
  wire [6:0] s_76;
  wire [0:0] s_77;
  wire [0:0] s_78;
  wire [5:0] s_79;
  wire [0:0] s_80;
  wire [0:0] s_81;
  wire [4:0] s_82;
  wire [0:0] s_83;
  wire [0:0] s_84;
  wire [3:0] s_85;
  wire [0:0] s_86;
  wire [0:0] s_87;
  wire [2:0] s_88;
  wire [0:0] s_89;
  wire [0:0] s_90;
  wire [1:0] s_91;
  wire [0:0] s_92;
  wire [0:0] s_93;
  wire [0:0] s_94;
  wire [1:0] s_95;
  wire [3:0] s_96;
  wire [7:0] s_97;
  wire [15:0] s_98;
  wire [31:0] s_99;
  wire [63:0] s_100;
  wire [62:0] s_101;
  wire [61:0] s_102;
  wire [60:0] s_103;
  wire [59:0] s_104;
  wire [58:0] s_105;
  wire [57:0] s_106;
  wire [56:0] s_107;
  wire [55:0] s_108;
  wire [54:0] s_109;
  wire [53:0] s_110;
  wire [52:0] s_111;
  wire [51:0] s_112;
  wire [50:0] s_113;
  wire [49:0] s_114;
  wire [48:0] s_115;
  wire [0:0] s_116;
  wire [0:0] s_117;
  wire [0:0] s_118;
  wire [0:0] s_119;
  wire [0:0] s_120;
  wire [0:0] s_121;
  wire [0:0] s_122;
  wire [0:0] s_123;
  wire [0:0] s_124;
  wire [0:0] s_125;
  wire [0:0] s_126;
  wire [0:0] s_127;
  wire [0:0] s_128;
  wire [0:0] s_129;
  wire [0:0] s_130;
  wire [0:0] s_131;
  wire [0:0] s_132;
  wire [0:0] s_133;
  wire [0:0] s_134;
  wire [0:0] s_135;
  wire [0:0] s_136;
  wire [0:0] s_137;
  wire [0:0] s_138;
  wire [1:0] s_139;
  wire [0:0] s_140;
  wire [0:0] s_141;
  wire [0:0] s_142;
  wire [1:0] s_143;
  wire [0:0] s_144;
  wire [0:0] s_145;
  wire [0:0] s_146;
  wire [0:0] s_147;
  wire [0:0] s_148;
  wire [0:0] s_149;
  wire [1:0] s_150;
  wire [0:0] s_151;
  wire [0:0] s_152;
  wire [0:0] s_153;
  wire [0:0] s_154;
  wire [0:0] s_155;
  wire [0:0] s_156;
  wire [2:0] s_157;
  wire [0:0] s_158;
  wire [0:0] s_159;
  wire [1:0] s_160;
  wire [0:0] s_161;
  wire [0:0] s_162;
  wire [0:0] s_163;
  wire [1:0] s_164;
  wire [3:0] s_165;
  wire [0:0] s_166;
  wire [0:0] s_167;
  wire [0:0] s_168;
  wire [0:0] s_169;
  wire [0:0] s_170;
  wire [0:0] s_171;
  wire [0:0] s_172;
  wire [1:0] s_173;
  wire [0:0] s_174;
  wire [0:0] s_175;
  wire [0:0] s_176;
  wire [1:0] s_177;
  wire [0:0] s_178;
  wire [0:0] s_179;
  wire [0:0] s_180;
  wire [0:0] s_181;
  wire [0:0] s_182;
  wire [0:0] s_183;
  wire [1:0] s_184;
  wire [0:0] s_185;
  wire [0:0] s_186;
  wire [0:0] s_187;
  wire [0:0] s_188;
  wire [0:0] s_189;
  wire [2:0] s_190;
  wire [0:0] s_191;
  wire [0:0] s_192;
  wire [1:0] s_193;
  wire [1:0] s_194;
  wire [1:0] s_195;
  wire [0:0] s_196;
  wire [3:0] s_197;
  wire [0:0] s_198;
  wire [0:0] s_199;
  wire [2:0] s_200;
  wire [0:0] s_201;
  wire [0:0] s_202;
  wire [1:0] s_203;
  wire [0:0] s_204;
  wire [0:0] s_205;
  wire [0:0] s_206;
  wire [1:0] s_207;
  wire [3:0] s_208;
  wire [7:0] s_209;
  wire [0:0] s_210;
  wire [0:0] s_211;
  wire [0:0] s_212;
  wire [0:0] s_213;
  wire [0:0] s_214;
  wire [0:0] s_215;
  wire [0:0] s_216;
  wire [1:0] s_217;
  wire [0:0] s_218;
  wire [0:0] s_219;
  wire [0:0] s_220;
  wire [1:0] s_221;
  wire [0:0] s_222;
  wire [0:0] s_223;
  wire [0:0] s_224;
  wire [0:0] s_225;
  wire [0:0] s_226;
  wire [0:0] s_227;
  wire [1:0] s_228;
  wire [0:0] s_229;
  wire [0:0] s_230;
  wire [0:0] s_231;
  wire [0:0] s_232;
  wire [0:0] s_233;
  wire [0:0] s_234;
  wire [2:0] s_235;
  wire [0:0] s_236;
  wire [0:0] s_237;
  wire [1:0] s_238;
  wire [0:0] s_239;
  wire [0:0] s_240;
  wire [0:0] s_241;
  wire [1:0] s_242;
  wire [3:0] s_243;
  wire [0:0] s_244;
  wire [0:0] s_245;
  wire [0:0] s_246;
  wire [0:0] s_247;
  wire [0:0] s_248;
  wire [0:0] s_249;
  wire [0:0] s_250;
  wire [1:0] s_251;
  wire [0:0] s_252;
  wire [0:0] s_253;
  wire [0:0] s_254;
  wire [1:0] s_255;
  wire [0:0] s_256;
  wire [0:0] s_257;
  wire [0:0] s_258;
  wire [0:0] s_259;
  wire [0:0] s_260;
  wire [0:0] s_261;
  wire [1:0] s_262;
  wire [0:0] s_263;
  wire [0:0] s_264;
  wire [0:0] s_265;
  wire [0:0] s_266;
  wire [0:0] s_267;
  wire [2:0] s_268;
  wire [0:0] s_269;
  wire [0:0] s_270;
  wire [1:0] s_271;
  wire [1:0] s_272;
  wire [1:0] s_273;
  wire [3:0] s_274;
  wire [0:0] s_275;
  wire [0:0] s_276;
  wire [2:0] s_277;
  wire [2:0] s_278;
  wire [2:0] s_279;
  wire [0:0] s_280;
  wire [4:0] s_281;
  wire [0:0] s_282;
  wire [0:0] s_283;
  wire [3:0] s_284;
  wire [0:0] s_285;
  wire [0:0] s_286;
  wire [2:0] s_287;
  wire [0:0] s_288;
  wire [0:0] s_289;
  wire [1:0] s_290;
  wire [0:0] s_291;
  wire [0:0] s_292;
  wire [0:0] s_293;
  wire [1:0] s_294;
  wire [3:0] s_295;
  wire [7:0] s_296;
  wire [15:0] s_297;
  wire [0:0] s_298;
  wire [0:0] s_299;
  wire [0:0] s_300;
  wire [0:0] s_301;
  wire [0:0] s_302;
  wire [0:0] s_303;
  wire [0:0] s_304;
  wire [1:0] s_305;
  wire [0:0] s_306;
  wire [0:0] s_307;
  wire [0:0] s_308;
  wire [1:0] s_309;
  wire [0:0] s_310;
  wire [0:0] s_311;
  wire [0:0] s_312;
  wire [0:0] s_313;
  wire [0:0] s_314;
  wire [0:0] s_315;
  wire [1:0] s_316;
  wire [0:0] s_317;
  wire [0:0] s_318;
  wire [0:0] s_319;
  wire [0:0] s_320;
  wire [0:0] s_321;
  wire [0:0] s_322;
  wire [2:0] s_323;
  wire [0:0] s_324;
  wire [0:0] s_325;
  wire [1:0] s_326;
  wire [0:0] s_327;
  wire [0:0] s_328;
  wire [0:0] s_329;
  wire [1:0] s_330;
  wire [3:0] s_331;
  wire [0:0] s_332;
  wire [0:0] s_333;
  wire [0:0] s_334;
  wire [0:0] s_335;
  wire [0:0] s_336;
  wire [0:0] s_337;
  wire [0:0] s_338;
  wire [1:0] s_339;
  wire [0:0] s_340;
  wire [0:0] s_341;
  wire [0:0] s_342;
  wire [1:0] s_343;
  wire [0:0] s_344;
  wire [0:0] s_345;
  wire [0:0] s_346;
  wire [0:0] s_347;
  wire [0:0] s_348;
  wire [0:0] s_349;
  wire [1:0] s_350;
  wire [0:0] s_351;
  wire [0:0] s_352;
  wire [0:0] s_353;
  wire [0:0] s_354;
  wire [0:0] s_355;
  wire [2:0] s_356;
  wire [0:0] s_357;
  wire [0:0] s_358;
  wire [1:0] s_359;
  wire [1:0] s_360;
  wire [1:0] s_361;
  wire [0:0] s_362;
  wire [3:0] s_363;
  wire [0:0] s_364;
  wire [0:0] s_365;
  wire [2:0] s_366;
  wire [0:0] s_367;
  wire [0:0] s_368;
  wire [1:0] s_369;
  wire [0:0] s_370;
  wire [0:0] s_371;
  wire [0:0] s_372;
  wire [1:0] s_373;
  wire [3:0] s_374;
  wire [7:0] s_375;
  wire [0:0] s_376;
  wire [0:0] s_377;
  wire [0:0] s_378;
  wire [0:0] s_379;
  wire [0:0] s_380;
  wire [0:0] s_381;
  wire [0:0] s_382;
  wire [1:0] s_383;
  wire [0:0] s_384;
  wire [0:0] s_385;
  wire [0:0] s_386;
  wire [1:0] s_387;
  wire [0:0] s_388;
  wire [0:0] s_389;
  wire [0:0] s_390;
  wire [0:0] s_391;
  wire [0:0] s_392;
  wire [0:0] s_393;
  wire [1:0] s_394;
  wire [0:0] s_395;
  wire [0:0] s_396;
  wire [0:0] s_397;
  wire [0:0] s_398;
  wire [0:0] s_399;
  wire [0:0] s_400;
  wire [2:0] s_401;
  wire [0:0] s_402;
  wire [0:0] s_403;
  wire [1:0] s_404;
  wire [0:0] s_405;
  wire [0:0] s_406;
  wire [0:0] s_407;
  wire [1:0] s_408;
  wire [3:0] s_409;
  wire [0:0] s_410;
  wire [0:0] s_411;
  wire [0:0] s_412;
  wire [0:0] s_413;
  wire [0:0] s_414;
  wire [0:0] s_415;
  wire [0:0] s_416;
  wire [1:0] s_417;
  wire [0:0] s_418;
  wire [0:0] s_419;
  wire [0:0] s_420;
  wire [1:0] s_421;
  wire [0:0] s_422;
  wire [0:0] s_423;
  wire [0:0] s_424;
  wire [0:0] s_425;
  wire [0:0] s_426;
  wire [0:0] s_427;
  wire [1:0] s_428;
  wire [0:0] s_429;
  wire [0:0] s_430;
  wire [0:0] s_431;
  wire [0:0] s_432;
  wire [0:0] s_433;
  wire [2:0] s_434;
  wire [0:0] s_435;
  wire [0:0] s_436;
  wire [1:0] s_437;
  wire [1:0] s_438;
  wire [1:0] s_439;
  wire [3:0] s_440;
  wire [0:0] s_441;
  wire [0:0] s_442;
  wire [2:0] s_443;
  wire [2:0] s_444;
  wire [2:0] s_445;
  wire [4:0] s_446;
  wire [0:0] s_447;
  wire [0:0] s_448;
  wire [3:0] s_449;
  wire [3:0] s_450;
  wire [3:0] s_451;
  wire [0:0] s_452;
  wire [5:0] s_453;
  wire [0:0] s_454;
  wire [0:0] s_455;
  wire [4:0] s_456;
  wire [0:0] s_457;
  wire [0:0] s_458;
  wire [3:0] s_459;
  wire [0:0] s_460;
  wire [0:0] s_461;
  wire [2:0] s_462;
  wire [0:0] s_463;
  wire [0:0] s_464;
  wire [1:0] s_465;
  wire [0:0] s_466;
  wire [0:0] s_467;
  wire [0:0] s_468;
  wire [1:0] s_469;
  wire [3:0] s_470;
  wire [7:0] s_471;
  wire [15:0] s_472;
  wire [31:0] s_473;
  wire [0:0] s_474;
  wire [0:0] s_475;
  wire [0:0] s_476;
  wire [0:0] s_477;
  wire [0:0] s_478;
  wire [0:0] s_479;
  wire [0:0] s_480;
  wire [1:0] s_481;
  wire [0:0] s_482;
  wire [0:0] s_483;
  wire [0:0] s_484;
  wire [1:0] s_485;
  wire [0:0] s_486;
  wire [0:0] s_487;
  wire [0:0] s_488;
  wire [0:0] s_489;
  wire [0:0] s_490;
  wire [0:0] s_491;
  wire [1:0] s_492;
  wire [0:0] s_493;
  wire [0:0] s_494;
  wire [0:0] s_495;
  wire [0:0] s_496;
  wire [0:0] s_497;
  wire [0:0] s_498;
  wire [2:0] s_499;
  wire [0:0] s_500;
  wire [0:0] s_501;
  wire [1:0] s_502;
  wire [0:0] s_503;
  wire [0:0] s_504;
  wire [0:0] s_505;
  wire [1:0] s_506;
  wire [3:0] s_507;
  wire [0:0] s_508;
  wire [0:0] s_509;
  wire [0:0] s_510;
  wire [0:0] s_511;
  wire [0:0] s_512;
  wire [0:0] s_513;
  wire [0:0] s_514;
  wire [1:0] s_515;
  wire [0:0] s_516;
  wire [0:0] s_517;
  wire [0:0] s_518;
  wire [1:0] s_519;
  wire [0:0] s_520;
  wire [0:0] s_521;
  wire [0:0] s_522;
  wire [0:0] s_523;
  wire [0:0] s_524;
  wire [0:0] s_525;
  wire [1:0] s_526;
  wire [0:0] s_527;
  wire [0:0] s_528;
  wire [0:0] s_529;
  wire [0:0] s_530;
  wire [0:0] s_531;
  wire [2:0] s_532;
  wire [0:0] s_533;
  wire [0:0] s_534;
  wire [1:0] s_535;
  wire [1:0] s_536;
  wire [1:0] s_537;
  wire [0:0] s_538;
  wire [3:0] s_539;
  wire [0:0] s_540;
  wire [0:0] s_541;
  wire [2:0] s_542;
  wire [0:0] s_543;
  wire [0:0] s_544;
  wire [1:0] s_545;
  wire [0:0] s_546;
  wire [0:0] s_547;
  wire [0:0] s_548;
  wire [1:0] s_549;
  wire [3:0] s_550;
  wire [7:0] s_551;
  wire [0:0] s_552;
  wire [0:0] s_553;
  wire [0:0] s_554;
  wire [0:0] s_555;
  wire [0:0] s_556;
  wire [0:0] s_557;
  wire [0:0] s_558;
  wire [1:0] s_559;
  wire [0:0] s_560;
  wire [0:0] s_561;
  wire [0:0] s_562;
  wire [1:0] s_563;
  wire [0:0] s_564;
  wire [0:0] s_565;
  wire [0:0] s_566;
  wire [0:0] s_567;
  wire [0:0] s_568;
  wire [0:0] s_569;
  wire [1:0] s_570;
  wire [0:0] s_571;
  wire [0:0] s_572;
  wire [0:0] s_573;
  wire [0:0] s_574;
  wire [0:0] s_575;
  wire [0:0] s_576;
  wire [2:0] s_577;
  wire [0:0] s_578;
  wire [0:0] s_579;
  wire [1:0] s_580;
  wire [0:0] s_581;
  wire [0:0] s_582;
  wire [0:0] s_583;
  wire [1:0] s_584;
  wire [3:0] s_585;
  wire [0:0] s_586;
  wire [0:0] s_587;
  wire [0:0] s_588;
  wire [0:0] s_589;
  wire [0:0] s_590;
  wire [0:0] s_591;
  wire [0:0] s_592;
  wire [1:0] s_593;
  wire [0:0] s_594;
  wire [0:0] s_595;
  wire [0:0] s_596;
  wire [1:0] s_597;
  wire [0:0] s_598;
  wire [0:0] s_599;
  wire [0:0] s_600;
  wire [0:0] s_601;
  wire [0:0] s_602;
  wire [0:0] s_603;
  wire [1:0] s_604;
  wire [0:0] s_605;
  wire [0:0] s_606;
  wire [0:0] s_607;
  wire [0:0] s_608;
  wire [0:0] s_609;
  wire [2:0] s_610;
  wire [0:0] s_611;
  wire [0:0] s_612;
  wire [1:0] s_613;
  wire [1:0] s_614;
  wire [1:0] s_615;
  wire [3:0] s_616;
  wire [0:0] s_617;
  wire [0:0] s_618;
  wire [2:0] s_619;
  wire [2:0] s_620;
  wire [2:0] s_621;
  wire [0:0] s_622;
  wire [4:0] s_623;
  wire [0:0] s_624;
  wire [0:0] s_625;
  wire [3:0] s_626;
  wire [0:0] s_627;
  wire [0:0] s_628;
  wire [2:0] s_629;
  wire [0:0] s_630;
  wire [0:0] s_631;
  wire [1:0] s_632;
  wire [0:0] s_633;
  wire [0:0] s_634;
  wire [0:0] s_635;
  wire [1:0] s_636;
  wire [3:0] s_637;
  wire [7:0] s_638;
  wire [15:0] s_639;
  wire [0:0] s_640;
  wire [0:0] s_641;
  wire [0:0] s_642;
  wire [0:0] s_643;
  wire [0:0] s_644;
  wire [0:0] s_645;
  wire [0:0] s_646;
  wire [1:0] s_647;
  wire [0:0] s_648;
  wire [0:0] s_649;
  wire [0:0] s_650;
  wire [1:0] s_651;
  wire [0:0] s_652;
  wire [0:0] s_653;
  wire [0:0] s_654;
  wire [0:0] s_655;
  wire [0:0] s_656;
  wire [0:0] s_657;
  wire [1:0] s_658;
  wire [0:0] s_659;
  wire [0:0] s_660;
  wire [0:0] s_661;
  wire [0:0] s_662;
  wire [0:0] s_663;
  wire [0:0] s_664;
  wire [2:0] s_665;
  wire [0:0] s_666;
  wire [0:0] s_667;
  wire [1:0] s_668;
  wire [0:0] s_669;
  wire [0:0] s_670;
  wire [0:0] s_671;
  wire [1:0] s_672;
  wire [3:0] s_673;
  wire [0:0] s_674;
  wire [0:0] s_675;
  wire [0:0] s_676;
  wire [0:0] s_677;
  wire [0:0] s_678;
  wire [0:0] s_679;
  wire [0:0] s_680;
  wire [1:0] s_681;
  wire [0:0] s_682;
  wire [0:0] s_683;
  wire [0:0] s_684;
  wire [1:0] s_685;
  wire [0:0] s_686;
  wire [0:0] s_687;
  wire [0:0] s_688;
  wire [0:0] s_689;
  wire [0:0] s_690;
  wire [0:0] s_691;
  wire [1:0] s_692;
  wire [0:0] s_693;
  wire [0:0] s_694;
  wire [0:0] s_695;
  wire [0:0] s_696;
  wire [0:0] s_697;
  wire [2:0] s_698;
  wire [0:0] s_699;
  wire [0:0] s_700;
  wire [1:0] s_701;
  wire [1:0] s_702;
  wire [1:0] s_703;
  wire [0:0] s_704;
  wire [3:0] s_705;
  wire [0:0] s_706;
  wire [0:0] s_707;
  wire [2:0] s_708;
  wire [0:0] s_709;
  wire [0:0] s_710;
  wire [1:0] s_711;
  wire [0:0] s_712;
  wire [0:0] s_713;
  wire [0:0] s_714;
  wire [1:0] s_715;
  wire [3:0] s_716;
  wire [7:0] s_717;
  wire [0:0] s_718;
  wire [0:0] s_719;
  wire [0:0] s_720;
  wire [0:0] s_721;
  wire [0:0] s_722;
  wire [0:0] s_723;
  wire [0:0] s_724;
  wire [1:0] s_725;
  wire [0:0] s_726;
  wire [0:0] s_727;
  wire [0:0] s_728;
  wire [1:0] s_729;
  wire [0:0] s_730;
  wire [0:0] s_731;
  wire [0:0] s_732;
  wire [0:0] s_733;
  wire [0:0] s_734;
  wire [0:0] s_735;
  wire [1:0] s_736;
  wire [0:0] s_737;
  wire [0:0] s_738;
  wire [0:0] s_739;
  wire [0:0] s_740;
  wire [0:0] s_741;
  wire [0:0] s_742;
  wire [2:0] s_743;
  wire [0:0] s_744;
  wire [0:0] s_745;
  wire [1:0] s_746;
  wire [0:0] s_747;
  wire [0:0] s_748;
  wire [0:0] s_749;
  wire [1:0] s_750;
  wire [3:0] s_751;
  wire [0:0] s_752;
  wire [0:0] s_753;
  wire [0:0] s_754;
  wire [0:0] s_755;
  wire [0:0] s_756;
  wire [0:0] s_757;
  wire [0:0] s_758;
  wire [1:0] s_759;
  wire [0:0] s_760;
  wire [0:0] s_761;
  wire [0:0] s_762;
  wire [1:0] s_763;
  wire [0:0] s_764;
  wire [0:0] s_765;
  wire [0:0] s_766;
  wire [0:0] s_767;
  wire [0:0] s_768;
  wire [0:0] s_769;
  wire [1:0] s_770;
  wire [0:0] s_771;
  wire [0:0] s_772;
  wire [0:0] s_773;
  wire [0:0] s_774;
  wire [0:0] s_775;
  wire [2:0] s_776;
  wire [0:0] s_777;
  wire [0:0] s_778;
  wire [1:0] s_779;
  wire [1:0] s_780;
  wire [1:0] s_781;
  wire [3:0] s_782;
  wire [0:0] s_783;
  wire [0:0] s_784;
  wire [2:0] s_785;
  wire [2:0] s_786;
  wire [2:0] s_787;
  wire [4:0] s_788;
  wire [0:0] s_789;
  wire [0:0] s_790;
  wire [3:0] s_791;
  wire [3:0] s_792;
  wire [3:0] s_793;
  wire [5:0] s_794;
  wire [0:0] s_795;
  wire [0:0] s_796;
  wire [4:0] s_797;
  wire [4:0] s_798;
  wire [4:0] s_799;
  wire [9:0] s_800;
  wire [9:0] s_801;
  wire [9:0] s_802;
  wire [9:0] s_803;
  wire [9:0] s_804;
  wire [0:0] s_805;
  wire [9:0] s_806;
  wire [9:0] s_807;
  wire [0:0] s_808;
  wire [23:0] s_809;
  wire [0:0] s_810;
  wire [0:0] s_811;
  wire [0:0] s_812;
  wire [0:0] s_813;
  wire [0:0] s_814;
  wire [0:0] s_815;
  wire [0:0] s_816;
  wire [0:0] s_817;
  wire [0:0] s_818;
  wire [21:0] s_819;
  wire [23:0] s_820;
  wire [0:0] s_821;
  wire [0:0] s_822;
  wire [23:0] s_823;
  wire [0:0] s_824;
  wire [31:0] s_825;
  wire [8:0] s_826;
  wire [0:0] s_827;
  wire [7:0] s_828;
  wire [7:0] s_829;
  wire [9:0] s_830;
  wire [9:0] s_831;
  wire [9:0] s_832;
  wire [9:0] s_833;
  wire [9:0] s_834;
  wire [9:0] s_835;
  wire [6:0] s_836;
  wire [22:0] s_837;
  wire [0:0] s_838;
  wire [0:0] s_839;
  wire [7:0] s_840;
  wire [0:0] s_841;
  wire [0:0] s_842;
  wire [0:0] s_843;
  wire [23:0] s_844;
  wire [0:0] s_845;
  wire [0:0] s_846;
  wire [0:0] s_847;
  wire [8:0] s_848;
  wire [0:0] s_849;
  wire [0:0] s_850;
  wire [0:0] s_851;
  wire [7:0] s_852;
  wire [0:0] s_853;
  wire [22:0] s_854;
  wire [0:0] s_855;
  wire [0:0] s_856;
  wire [0:0] s_857;
  wire [7:0] s_858;
  wire [0:0] s_859;
  wire [22:0] s_860;
  wire [0:0] s_861;
  wire [0:0] s_862;
  wire [0:0] s_863;
  wire [0:0] s_864;
  wire [7:0] s_865;
  wire [0:0] s_866;
  wire [22:0] s_867;
  wire [0:0] s_868;
  wire [0:0] s_869;
  wire [7:0] s_870;
  wire [0:0] s_871;
  wire [22:0] s_872;

  assign s_0 = s_861?s_1:s_9;
  dq #(32, 6) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_8};
  assign s_3 = s_4 ^ s_6;
  assign s_4 = s_5[31];
  assign s_5 = mul_a;
  assign s_6 = s_7[31];
  assign s_7 = mul_b;
  assign s_8 = 31'd2143289344;
  assign s_9 = s_845?s_10:s_13;
  dq #(32, 6) dq_s_10 (clk, s_10, s_11);
  assign s_11 = {s_3,s_12};
  assign s_12 = 31'd2139095040;
  assign s_13 = s_843?s_14:s_17;
  dq #(32, 6) dq_s_14 (clk, s_14, s_15);
  assign s_15 = {s_3,s_16};
  assign s_16 = 31'd0;
  assign s_17 = s_838?s_18:s_825;
  assign s_18 = {s_19,s_22};
  dq #(9, 6) dq_s_19 (clk, s_19, s_20);
  assign s_20 = {s_3,s_21};
  assign s_21 = 8'd0;
  assign s_22 = s_23[22:0];
  dq #(24, 1) dq_s_23 (clk, s_23, s_24);
  assign s_24 = s_824?s_25:s_823;
  assign s_25 = s_26[24:1];
  assign s_26 = s_810?s_27:s_809;
  dq #(25, 1) dq_s_27 (clk, s_27, s_28);
  assign s_28 = s_29 + s_808;
  assign s_29 = s_30;
  assign s_30 = s_31[47:24];
  dq #(48, 1) dq_s_31 (clk, s_31, s_32);
  assign s_32 = s_33 << s_73;
  dq #(48, 2) dq_s_33 (clk, s_33, s_34);
  dq #(48, 1) dq_s_34 (clk, s_34, s_35);
  assign s_35 = s_36 >> s_59;
  assign s_36 = s_37 * s_48;
  assign s_37 = s_38;
  assign s_38 = {s_39,s_47};
  assign s_39 = s_42?s_40:s_41;
  assign s_40 = 1'd0;
  assign s_41 = 1'd1;
  assign s_42 = s_43 == s_46;
  assign s_43 = s_44 - s_45;
  assign s_44 = s_5[30:23];
  assign s_45 = 7'd127;
  assign s_46 = -8'd127;
  assign s_47 = s_5[22:0];
  assign s_48 = s_49;
  assign s_49 = {s_50,s_58};
  assign s_50 = s_53?s_51:s_52;
  assign s_51 = 1'd0;
  assign s_52 = 1'd1;
  assign s_53 = s_54 == s_57;
  assign s_54 = s_55 - s_56;
  assign s_55 = s_7[30:23];
  assign s_56 = 7'd127;
  assign s_57 = -8'd127;
  assign s_58 = s_7[22:0];
  assign s_59 = s_72?s_60:s_61;
  assign s_60 = 1'd0;
  assign s_61 = s_62 - s_63;
  assign s_62 = -10'd126;
  assign s_63 = s_64 + s_71;
  assign s_64 = s_65 + s_68;
  assign s_65 = $signed(s_66);
  assign s_66 = s_42?s_67:s_43;
  assign s_67 = -8'd126;
  assign s_68 = $signed(s_69);
  assign s_69 = s_53?s_70:s_54;
  assign s_70 = -8'd126;
  assign s_71 = 1'd1;
  assign s_72 = s_61[9];
  dq #(10, 1) dq_s_73 (clk, s_73, s_74);
  assign s_74 = s_805?s_75:s_800;
  dq #(7, 1) dq_s_75 (clk, s_75, s_76);
  assign s_76 = {s_77,s_794};
  assign s_77 = s_78 & s_452;
  assign s_78 = s_79[5];
  assign s_79 = {s_80,s_446};
  assign s_80 = s_81 & s_280;
  assign s_81 = s_82[4];
  assign s_82 = {s_83,s_274};
  assign s_83 = s_84 & s_196;
  assign s_84 = s_85[3];
  assign s_85 = {s_86,s_190};
  assign s_86 = s_87 & s_156;
  assign s_87 = s_88[2];
  assign s_88 = {s_89,s_150};
  assign s_89 = s_90 & s_138;
  assign s_90 = s_91[1];
  assign s_91 = {s_92,s_134};
  assign s_92 = s_93 & s_132;
  assign s_93 = ~s_94;
  assign s_94 = s_95[1];
  assign s_95 = s_96[3:2];
  assign s_96 = s_97[7:4];
  assign s_97 = s_98[15:8];
  assign s_98 = s_99[31:16];
  assign s_99 = s_100[63:32];
  assign s_100 = {s_101,s_131};
  assign s_101 = {s_102,s_130};
  assign s_102 = {s_103,s_129};
  assign s_103 = {s_104,s_128};
  assign s_104 = {s_105,s_127};
  assign s_105 = {s_106,s_126};
  assign s_106 = {s_107,s_125};
  assign s_107 = {s_108,s_124};
  assign s_108 = {s_109,s_123};
  assign s_109 = {s_110,s_122};
  assign s_110 = {s_111,s_121};
  assign s_111 = {s_112,s_120};
  assign s_112 = {s_113,s_119};
  assign s_113 = {s_114,s_118};
  assign s_114 = {s_115,s_117};
  assign s_115 = {s_34,s_116};
  assign s_116 = 1'd1;
  assign s_117 = 1'd1;
  assign s_118 = 1'd1;
  assign s_119 = 1'd1;
  assign s_120 = 1'd1;
  assign s_121 = 1'd1;
  assign s_122 = 1'd1;
  assign s_123 = 1'd1;
  assign s_124 = 1'd1;
  assign s_125 = 1'd1;
  assign s_126 = 1'd1;
  assign s_127 = 1'd1;
  assign s_128 = 1'd1;
  assign s_129 = 1'd1;
  assign s_130 = 1'd1;
  assign s_131 = 1'd1;
  assign s_132 = ~s_133;
  assign s_133 = s_95[0];
  assign s_134 = s_135 & s_137;
  assign s_135 = ~s_136;
  assign s_136 = s_95[1];
  assign s_137 = s_95[0];
  assign s_138 = s_139[1];
  assign s_139 = {s_140,s_146};
  assign s_140 = s_141 & s_144;
  assign s_141 = ~s_142;
  assign s_142 = s_143[1];
  assign s_143 = s_96[1:0];
  assign s_144 = ~s_145;
  assign s_145 = s_143[0];
  assign s_146 = s_147 & s_149;
  assign s_147 = ~s_148;
  assign s_148 = s_143[1];
  assign s_149 = s_143[0];
  assign s_150 = {s_151,s_153};
  assign s_151 = s_90 & s_152;
  assign s_152 = ~s_138;
  assign s_153 = s_90?s_154:s_155;
  assign s_154 = s_139[0:0];
  assign s_155 = s_91[0:0];
  assign s_156 = s_157[2];
  assign s_157 = {s_158,s_184};
  assign s_158 = s_159 & s_172;
  assign s_159 = s_160[1];
  assign s_160 = {s_161,s_168};
  assign s_161 = s_162 & s_166;
  assign s_162 = ~s_163;
  assign s_163 = s_164[1];
  assign s_164 = s_165[3:2];
  assign s_165 = s_97[3:0];
  assign s_166 = ~s_167;
  assign s_167 = s_164[0];
  assign s_168 = s_169 & s_171;
  assign s_169 = ~s_170;
  assign s_170 = s_164[1];
  assign s_171 = s_164[0];
  assign s_172 = s_173[1];
  assign s_173 = {s_174,s_180};
  assign s_174 = s_175 & s_178;
  assign s_175 = ~s_176;
  assign s_176 = s_177[1];
  assign s_177 = s_165[1:0];
  assign s_178 = ~s_179;
  assign s_179 = s_177[0];
  assign s_180 = s_181 & s_183;
  assign s_181 = ~s_182;
  assign s_182 = s_177[1];
  assign s_183 = s_177[0];
  assign s_184 = {s_185,s_187};
  assign s_185 = s_159 & s_186;
  assign s_186 = ~s_172;
  assign s_187 = s_159?s_188:s_189;
  assign s_188 = s_173[0:0];
  assign s_189 = s_160[0:0];
  assign s_190 = {s_191,s_193};
  assign s_191 = s_87 & s_192;
  assign s_192 = ~s_156;
  assign s_193 = s_87?s_194:s_195;
  assign s_194 = s_157[1:0];
  assign s_195 = s_88[1:0];
  assign s_196 = s_197[3];
  assign s_197 = {s_198,s_268};
  assign s_198 = s_199 & s_234;
  assign s_199 = s_200[2];
  assign s_200 = {s_201,s_228};
  assign s_201 = s_202 & s_216;
  assign s_202 = s_203[1];
  assign s_203 = {s_204,s_212};
  assign s_204 = s_205 & s_210;
  assign s_205 = ~s_206;
  assign s_206 = s_207[1];
  assign s_207 = s_208[3:2];
  assign s_208 = s_209[7:4];
  assign s_209 = s_98[7:0];
  assign s_210 = ~s_211;
  assign s_211 = s_207[0];
  assign s_212 = s_213 & s_215;
  assign s_213 = ~s_214;
  assign s_214 = s_207[1];
  assign s_215 = s_207[0];
  assign s_216 = s_217[1];
  assign s_217 = {s_218,s_224};
  assign s_218 = s_219 & s_222;
  assign s_219 = ~s_220;
  assign s_220 = s_221[1];
  assign s_221 = s_208[1:0];
  assign s_222 = ~s_223;
  assign s_223 = s_221[0];
  assign s_224 = s_225 & s_227;
  assign s_225 = ~s_226;
  assign s_226 = s_221[1];
  assign s_227 = s_221[0];
  assign s_228 = {s_229,s_231};
  assign s_229 = s_202 & s_230;
  assign s_230 = ~s_216;
  assign s_231 = s_202?s_232:s_233;
  assign s_232 = s_217[0:0];
  assign s_233 = s_203[0:0];
  assign s_234 = s_235[2];
  assign s_235 = {s_236,s_262};
  assign s_236 = s_237 & s_250;
  assign s_237 = s_238[1];
  assign s_238 = {s_239,s_246};
  assign s_239 = s_240 & s_244;
  assign s_240 = ~s_241;
  assign s_241 = s_242[1];
  assign s_242 = s_243[3:2];
  assign s_243 = s_209[3:0];
  assign s_244 = ~s_245;
  assign s_245 = s_242[0];
  assign s_246 = s_247 & s_249;
  assign s_247 = ~s_248;
  assign s_248 = s_242[1];
  assign s_249 = s_242[0];
  assign s_250 = s_251[1];
  assign s_251 = {s_252,s_258};
  assign s_252 = s_253 & s_256;
  assign s_253 = ~s_254;
  assign s_254 = s_255[1];
  assign s_255 = s_243[1:0];
  assign s_256 = ~s_257;
  assign s_257 = s_255[0];
  assign s_258 = s_259 & s_261;
  assign s_259 = ~s_260;
  assign s_260 = s_255[1];
  assign s_261 = s_255[0];
  assign s_262 = {s_263,s_265};
  assign s_263 = s_237 & s_264;
  assign s_264 = ~s_250;
  assign s_265 = s_237?s_266:s_267;
  assign s_266 = s_251[0:0];
  assign s_267 = s_238[0:0];
  assign s_268 = {s_269,s_271};
  assign s_269 = s_199 & s_270;
  assign s_270 = ~s_234;
  assign s_271 = s_199?s_272:s_273;
  assign s_272 = s_235[1:0];
  assign s_273 = s_200[1:0];
  assign s_274 = {s_275,s_277};
  assign s_275 = s_84 & s_276;
  assign s_276 = ~s_196;
  assign s_277 = s_84?s_278:s_279;
  assign s_278 = s_197[2:0];
  assign s_279 = s_85[2:0];
  assign s_280 = s_281[4];
  assign s_281 = {s_282,s_440};
  assign s_282 = s_283 & s_362;
  assign s_283 = s_284[3];
  assign s_284 = {s_285,s_356};
  assign s_285 = s_286 & s_322;
  assign s_286 = s_287[2];
  assign s_287 = {s_288,s_316};
  assign s_288 = s_289 & s_304;
  assign s_289 = s_290[1];
  assign s_290 = {s_291,s_300};
  assign s_291 = s_292 & s_298;
  assign s_292 = ~s_293;
  assign s_293 = s_294[1];
  assign s_294 = s_295[3:2];
  assign s_295 = s_296[7:4];
  assign s_296 = s_297[15:8];
  assign s_297 = s_99[15:0];
  assign s_298 = ~s_299;
  assign s_299 = s_294[0];
  assign s_300 = s_301 & s_303;
  assign s_301 = ~s_302;
  assign s_302 = s_294[1];
  assign s_303 = s_294[0];
  assign s_304 = s_305[1];
  assign s_305 = {s_306,s_312};
  assign s_306 = s_307 & s_310;
  assign s_307 = ~s_308;
  assign s_308 = s_309[1];
  assign s_309 = s_295[1:0];
  assign s_310 = ~s_311;
  assign s_311 = s_309[0];
  assign s_312 = s_313 & s_315;
  assign s_313 = ~s_314;
  assign s_314 = s_309[1];
  assign s_315 = s_309[0];
  assign s_316 = {s_317,s_319};
  assign s_317 = s_289 & s_318;
  assign s_318 = ~s_304;
  assign s_319 = s_289?s_320:s_321;
  assign s_320 = s_305[0:0];
  assign s_321 = s_290[0:0];
  assign s_322 = s_323[2];
  assign s_323 = {s_324,s_350};
  assign s_324 = s_325 & s_338;
  assign s_325 = s_326[1];
  assign s_326 = {s_327,s_334};
  assign s_327 = s_328 & s_332;
  assign s_328 = ~s_329;
  assign s_329 = s_330[1];
  assign s_330 = s_331[3:2];
  assign s_331 = s_296[3:0];
  assign s_332 = ~s_333;
  assign s_333 = s_330[0];
  assign s_334 = s_335 & s_337;
  assign s_335 = ~s_336;
  assign s_336 = s_330[1];
  assign s_337 = s_330[0];
  assign s_338 = s_339[1];
  assign s_339 = {s_340,s_346};
  assign s_340 = s_341 & s_344;
  assign s_341 = ~s_342;
  assign s_342 = s_343[1];
  assign s_343 = s_331[1:0];
  assign s_344 = ~s_345;
  assign s_345 = s_343[0];
  assign s_346 = s_347 & s_349;
  assign s_347 = ~s_348;
  assign s_348 = s_343[1];
  assign s_349 = s_343[0];
  assign s_350 = {s_351,s_353};
  assign s_351 = s_325 & s_352;
  assign s_352 = ~s_338;
  assign s_353 = s_325?s_354:s_355;
  assign s_354 = s_339[0:0];
  assign s_355 = s_326[0:0];
  assign s_356 = {s_357,s_359};
  assign s_357 = s_286 & s_358;
  assign s_358 = ~s_322;
  assign s_359 = s_286?s_360:s_361;
  assign s_360 = s_323[1:0];
  assign s_361 = s_287[1:0];
  assign s_362 = s_363[3];
  assign s_363 = {s_364,s_434};
  assign s_364 = s_365 & s_400;
  assign s_365 = s_366[2];
  assign s_366 = {s_367,s_394};
  assign s_367 = s_368 & s_382;
  assign s_368 = s_369[1];
  assign s_369 = {s_370,s_378};
  assign s_370 = s_371 & s_376;
  assign s_371 = ~s_372;
  assign s_372 = s_373[1];
  assign s_373 = s_374[3:2];
  assign s_374 = s_375[7:4];
  assign s_375 = s_297[7:0];
  assign s_376 = ~s_377;
  assign s_377 = s_373[0];
  assign s_378 = s_379 & s_381;
  assign s_379 = ~s_380;
  assign s_380 = s_373[1];
  assign s_381 = s_373[0];
  assign s_382 = s_383[1];
  assign s_383 = {s_384,s_390};
  assign s_384 = s_385 & s_388;
  assign s_385 = ~s_386;
  assign s_386 = s_387[1];
  assign s_387 = s_374[1:0];
  assign s_388 = ~s_389;
  assign s_389 = s_387[0];
  assign s_390 = s_391 & s_393;
  assign s_391 = ~s_392;
  assign s_392 = s_387[1];
  assign s_393 = s_387[0];
  assign s_394 = {s_395,s_397};
  assign s_395 = s_368 & s_396;
  assign s_396 = ~s_382;
  assign s_397 = s_368?s_398:s_399;
  assign s_398 = s_383[0:0];
  assign s_399 = s_369[0:0];
  assign s_400 = s_401[2];
  assign s_401 = {s_402,s_428};
  assign s_402 = s_403 & s_416;
  assign s_403 = s_404[1];
  assign s_404 = {s_405,s_412};
  assign s_405 = s_406 & s_410;
  assign s_406 = ~s_407;
  assign s_407 = s_408[1];
  assign s_408 = s_409[3:2];
  assign s_409 = s_375[3:0];
  assign s_410 = ~s_411;
  assign s_411 = s_408[0];
  assign s_412 = s_413 & s_415;
  assign s_413 = ~s_414;
  assign s_414 = s_408[1];
  assign s_415 = s_408[0];
  assign s_416 = s_417[1];
  assign s_417 = {s_418,s_424};
  assign s_418 = s_419 & s_422;
  assign s_419 = ~s_420;
  assign s_420 = s_421[1];
  assign s_421 = s_409[1:0];
  assign s_422 = ~s_423;
  assign s_423 = s_421[0];
  assign s_424 = s_425 & s_427;
  assign s_425 = ~s_426;
  assign s_426 = s_421[1];
  assign s_427 = s_421[0];
  assign s_428 = {s_429,s_431};
  assign s_429 = s_403 & s_430;
  assign s_430 = ~s_416;
  assign s_431 = s_403?s_432:s_433;
  assign s_432 = s_417[0:0];
  assign s_433 = s_404[0:0];
  assign s_434 = {s_435,s_437};
  assign s_435 = s_365 & s_436;
  assign s_436 = ~s_400;
  assign s_437 = s_365?s_438:s_439;
  assign s_438 = s_401[1:0];
  assign s_439 = s_366[1:0];
  assign s_440 = {s_441,s_443};
  assign s_441 = s_283 & s_442;
  assign s_442 = ~s_362;
  assign s_443 = s_283?s_444:s_445;
  assign s_444 = s_363[2:0];
  assign s_445 = s_284[2:0];
  assign s_446 = {s_447,s_449};
  assign s_447 = s_81 & s_448;
  assign s_448 = ~s_280;
  assign s_449 = s_81?s_450:s_451;
  assign s_450 = s_281[3:0];
  assign s_451 = s_82[3:0];
  assign s_452 = s_453[5];
  assign s_453 = {s_454,s_788};
  assign s_454 = s_455 & s_622;
  assign s_455 = s_456[4];
  assign s_456 = {s_457,s_616};
  assign s_457 = s_458 & s_538;
  assign s_458 = s_459[3];
  assign s_459 = {s_460,s_532};
  assign s_460 = s_461 & s_498;
  assign s_461 = s_462[2];
  assign s_462 = {s_463,s_492};
  assign s_463 = s_464 & s_480;
  assign s_464 = s_465[1];
  assign s_465 = {s_466,s_476};
  assign s_466 = s_467 & s_474;
  assign s_467 = ~s_468;
  assign s_468 = s_469[1];
  assign s_469 = s_470[3:2];
  assign s_470 = s_471[7:4];
  assign s_471 = s_472[15:8];
  assign s_472 = s_473[31:16];
  assign s_473 = s_100[31:0];
  assign s_474 = ~s_475;
  assign s_475 = s_469[0];
  assign s_476 = s_477 & s_479;
  assign s_477 = ~s_478;
  assign s_478 = s_469[1];
  assign s_479 = s_469[0];
  assign s_480 = s_481[1];
  assign s_481 = {s_482,s_488};
  assign s_482 = s_483 & s_486;
  assign s_483 = ~s_484;
  assign s_484 = s_485[1];
  assign s_485 = s_470[1:0];
  assign s_486 = ~s_487;
  assign s_487 = s_485[0];
  assign s_488 = s_489 & s_491;
  assign s_489 = ~s_490;
  assign s_490 = s_485[1];
  assign s_491 = s_485[0];
  assign s_492 = {s_493,s_495};
  assign s_493 = s_464 & s_494;
  assign s_494 = ~s_480;
  assign s_495 = s_464?s_496:s_497;
  assign s_496 = s_481[0:0];
  assign s_497 = s_465[0:0];
  assign s_498 = s_499[2];
  assign s_499 = {s_500,s_526};
  assign s_500 = s_501 & s_514;
  assign s_501 = s_502[1];
  assign s_502 = {s_503,s_510};
  assign s_503 = s_504 & s_508;
  assign s_504 = ~s_505;
  assign s_505 = s_506[1];
  assign s_506 = s_507[3:2];
  assign s_507 = s_471[3:0];
  assign s_508 = ~s_509;
  assign s_509 = s_506[0];
  assign s_510 = s_511 & s_513;
  assign s_511 = ~s_512;
  assign s_512 = s_506[1];
  assign s_513 = s_506[0];
  assign s_514 = s_515[1];
  assign s_515 = {s_516,s_522};
  assign s_516 = s_517 & s_520;
  assign s_517 = ~s_518;
  assign s_518 = s_519[1];
  assign s_519 = s_507[1:0];
  assign s_520 = ~s_521;
  assign s_521 = s_519[0];
  assign s_522 = s_523 & s_525;
  assign s_523 = ~s_524;
  assign s_524 = s_519[1];
  assign s_525 = s_519[0];
  assign s_526 = {s_527,s_529};
  assign s_527 = s_501 & s_528;
  assign s_528 = ~s_514;
  assign s_529 = s_501?s_530:s_531;
  assign s_530 = s_515[0:0];
  assign s_531 = s_502[0:0];
  assign s_532 = {s_533,s_535};
  assign s_533 = s_461 & s_534;
  assign s_534 = ~s_498;
  assign s_535 = s_461?s_536:s_537;
  assign s_536 = s_499[1:0];
  assign s_537 = s_462[1:0];
  assign s_538 = s_539[3];
  assign s_539 = {s_540,s_610};
  assign s_540 = s_541 & s_576;
  assign s_541 = s_542[2];
  assign s_542 = {s_543,s_570};
  assign s_543 = s_544 & s_558;
  assign s_544 = s_545[1];
  assign s_545 = {s_546,s_554};
  assign s_546 = s_547 & s_552;
  assign s_547 = ~s_548;
  assign s_548 = s_549[1];
  assign s_549 = s_550[3:2];
  assign s_550 = s_551[7:4];
  assign s_551 = s_472[7:0];
  assign s_552 = ~s_553;
  assign s_553 = s_549[0];
  assign s_554 = s_555 & s_557;
  assign s_555 = ~s_556;
  assign s_556 = s_549[1];
  assign s_557 = s_549[0];
  assign s_558 = s_559[1];
  assign s_559 = {s_560,s_566};
  assign s_560 = s_561 & s_564;
  assign s_561 = ~s_562;
  assign s_562 = s_563[1];
  assign s_563 = s_550[1:0];
  assign s_564 = ~s_565;
  assign s_565 = s_563[0];
  assign s_566 = s_567 & s_569;
  assign s_567 = ~s_568;
  assign s_568 = s_563[1];
  assign s_569 = s_563[0];
  assign s_570 = {s_571,s_573};
  assign s_571 = s_544 & s_572;
  assign s_572 = ~s_558;
  assign s_573 = s_544?s_574:s_575;
  assign s_574 = s_559[0:0];
  assign s_575 = s_545[0:0];
  assign s_576 = s_577[2];
  assign s_577 = {s_578,s_604};
  assign s_578 = s_579 & s_592;
  assign s_579 = s_580[1];
  assign s_580 = {s_581,s_588};
  assign s_581 = s_582 & s_586;
  assign s_582 = ~s_583;
  assign s_583 = s_584[1];
  assign s_584 = s_585[3:2];
  assign s_585 = s_551[3:0];
  assign s_586 = ~s_587;
  assign s_587 = s_584[0];
  assign s_588 = s_589 & s_591;
  assign s_589 = ~s_590;
  assign s_590 = s_584[1];
  assign s_591 = s_584[0];
  assign s_592 = s_593[1];
  assign s_593 = {s_594,s_600};
  assign s_594 = s_595 & s_598;
  assign s_595 = ~s_596;
  assign s_596 = s_597[1];
  assign s_597 = s_585[1:0];
  assign s_598 = ~s_599;
  assign s_599 = s_597[0];
  assign s_600 = s_601 & s_603;
  assign s_601 = ~s_602;
  assign s_602 = s_597[1];
  assign s_603 = s_597[0];
  assign s_604 = {s_605,s_607};
  assign s_605 = s_579 & s_606;
  assign s_606 = ~s_592;
  assign s_607 = s_579?s_608:s_609;
  assign s_608 = s_593[0:0];
  assign s_609 = s_580[0:0];
  assign s_610 = {s_611,s_613};
  assign s_611 = s_541 & s_612;
  assign s_612 = ~s_576;
  assign s_613 = s_541?s_614:s_615;
  assign s_614 = s_577[1:0];
  assign s_615 = s_542[1:0];
  assign s_616 = {s_617,s_619};
  assign s_617 = s_458 & s_618;
  assign s_618 = ~s_538;
  assign s_619 = s_458?s_620:s_621;
  assign s_620 = s_539[2:0];
  assign s_621 = s_459[2:0];
  assign s_622 = s_623[4];
  assign s_623 = {s_624,s_782};
  assign s_624 = s_625 & s_704;
  assign s_625 = s_626[3];
  assign s_626 = {s_627,s_698};
  assign s_627 = s_628 & s_664;
  assign s_628 = s_629[2];
  assign s_629 = {s_630,s_658};
  assign s_630 = s_631 & s_646;
  assign s_631 = s_632[1];
  assign s_632 = {s_633,s_642};
  assign s_633 = s_634 & s_640;
  assign s_634 = ~s_635;
  assign s_635 = s_636[1];
  assign s_636 = s_637[3:2];
  assign s_637 = s_638[7:4];
  assign s_638 = s_639[15:8];
  assign s_639 = s_473[15:0];
  assign s_640 = ~s_641;
  assign s_641 = s_636[0];
  assign s_642 = s_643 & s_645;
  assign s_643 = ~s_644;
  assign s_644 = s_636[1];
  assign s_645 = s_636[0];
  assign s_646 = s_647[1];
  assign s_647 = {s_648,s_654};
  assign s_648 = s_649 & s_652;
  assign s_649 = ~s_650;
  assign s_650 = s_651[1];
  assign s_651 = s_637[1:0];
  assign s_652 = ~s_653;
  assign s_653 = s_651[0];
  assign s_654 = s_655 & s_657;
  assign s_655 = ~s_656;
  assign s_656 = s_651[1];
  assign s_657 = s_651[0];
  assign s_658 = {s_659,s_661};
  assign s_659 = s_631 & s_660;
  assign s_660 = ~s_646;
  assign s_661 = s_631?s_662:s_663;
  assign s_662 = s_647[0:0];
  assign s_663 = s_632[0:0];
  assign s_664 = s_665[2];
  assign s_665 = {s_666,s_692};
  assign s_666 = s_667 & s_680;
  assign s_667 = s_668[1];
  assign s_668 = {s_669,s_676};
  assign s_669 = s_670 & s_674;
  assign s_670 = ~s_671;
  assign s_671 = s_672[1];
  assign s_672 = s_673[3:2];
  assign s_673 = s_638[3:0];
  assign s_674 = ~s_675;
  assign s_675 = s_672[0];
  assign s_676 = s_677 & s_679;
  assign s_677 = ~s_678;
  assign s_678 = s_672[1];
  assign s_679 = s_672[0];
  assign s_680 = s_681[1];
  assign s_681 = {s_682,s_688};
  assign s_682 = s_683 & s_686;
  assign s_683 = ~s_684;
  assign s_684 = s_685[1];
  assign s_685 = s_673[1:0];
  assign s_686 = ~s_687;
  assign s_687 = s_685[0];
  assign s_688 = s_689 & s_691;
  assign s_689 = ~s_690;
  assign s_690 = s_685[1];
  assign s_691 = s_685[0];
  assign s_692 = {s_693,s_695};
  assign s_693 = s_667 & s_694;
  assign s_694 = ~s_680;
  assign s_695 = s_667?s_696:s_697;
  assign s_696 = s_681[0:0];
  assign s_697 = s_668[0:0];
  assign s_698 = {s_699,s_701};
  assign s_699 = s_628 & s_700;
  assign s_700 = ~s_664;
  assign s_701 = s_628?s_702:s_703;
  assign s_702 = s_665[1:0];
  assign s_703 = s_629[1:0];
  assign s_704 = s_705[3];
  assign s_705 = {s_706,s_776};
  assign s_706 = s_707 & s_742;
  assign s_707 = s_708[2];
  assign s_708 = {s_709,s_736};
  assign s_709 = s_710 & s_724;
  assign s_710 = s_711[1];
  assign s_711 = {s_712,s_720};
  assign s_712 = s_713 & s_718;
  assign s_713 = ~s_714;
  assign s_714 = s_715[1];
  assign s_715 = s_716[3:2];
  assign s_716 = s_717[7:4];
  assign s_717 = s_639[7:0];
  assign s_718 = ~s_719;
  assign s_719 = s_715[0];
  assign s_720 = s_721 & s_723;
  assign s_721 = ~s_722;
  assign s_722 = s_715[1];
  assign s_723 = s_715[0];
  assign s_724 = s_725[1];
  assign s_725 = {s_726,s_732};
  assign s_726 = s_727 & s_730;
  assign s_727 = ~s_728;
  assign s_728 = s_729[1];
  assign s_729 = s_716[1:0];
  assign s_730 = ~s_731;
  assign s_731 = s_729[0];
  assign s_732 = s_733 & s_735;
  assign s_733 = ~s_734;
  assign s_734 = s_729[1];
  assign s_735 = s_729[0];
  assign s_736 = {s_737,s_739};
  assign s_737 = s_710 & s_738;
  assign s_738 = ~s_724;
  assign s_739 = s_710?s_740:s_741;
  assign s_740 = s_725[0:0];
  assign s_741 = s_711[0:0];
  assign s_742 = s_743[2];
  assign s_743 = {s_744,s_770};
  assign s_744 = s_745 & s_758;
  assign s_745 = s_746[1];
  assign s_746 = {s_747,s_754};
  assign s_747 = s_748 & s_752;
  assign s_748 = ~s_749;
  assign s_749 = s_750[1];
  assign s_750 = s_751[3:2];
  assign s_751 = s_717[3:0];
  assign s_752 = ~s_753;
  assign s_753 = s_750[0];
  assign s_754 = s_755 & s_757;
  assign s_755 = ~s_756;
  assign s_756 = s_750[1];
  assign s_757 = s_750[0];
  assign s_758 = s_759[1];
  assign s_759 = {s_760,s_766};
  assign s_760 = s_761 & s_764;
  assign s_761 = ~s_762;
  assign s_762 = s_763[1];
  assign s_763 = s_751[1:0];
  assign s_764 = ~s_765;
  assign s_765 = s_763[0];
  assign s_766 = s_767 & s_769;
  assign s_767 = ~s_768;
  assign s_768 = s_763[1];
  assign s_769 = s_763[0];
  assign s_770 = {s_771,s_773};
  assign s_771 = s_745 & s_772;
  assign s_772 = ~s_758;
  assign s_773 = s_745?s_774:s_775;
  assign s_774 = s_759[0:0];
  assign s_775 = s_746[0:0];
  assign s_776 = {s_777,s_779};
  assign s_777 = s_707 & s_778;
  assign s_778 = ~s_742;
  assign s_779 = s_707?s_780:s_781;
  assign s_780 = s_743[1:0];
  assign s_781 = s_708[1:0];
  assign s_782 = {s_783,s_785};
  assign s_783 = s_625 & s_784;
  assign s_784 = ~s_704;
  assign s_785 = s_625?s_786:s_787;
  assign s_786 = s_705[2:0];
  assign s_787 = s_626[2:0];
  assign s_788 = {s_789,s_791};
  assign s_789 = s_455 & s_790;
  assign s_790 = ~s_622;
  assign s_791 = s_455?s_792:s_793;
  assign s_792 = s_623[3:0];
  assign s_793 = s_456[3:0];
  assign s_794 = {s_795,s_797};
  assign s_795 = s_78 & s_796;
  assign s_796 = ~s_452;
  assign s_797 = s_78?s_798:s_799;
  assign s_798 = s_453[4:0];
  assign s_799 = s_79[4:0];
  dq #(10, 1) dq_s_800 (clk, s_800, s_801);
  assign s_801 = s_802 - s_804;
  dq #(10, 1) dq_s_802 (clk, s_802, s_803);
  assign s_803 = s_63 + s_59;
  assign s_804 = -10'd126;
  assign s_805 = s_806 <= s_807;
  assign s_806 = s_75;
  dq #(10, 1) dq_s_807 (clk, s_807, s_801);
  assign s_808 = 1'd1;
  dq #(24, 1) dq_s_809 (clk, s_809, s_30);
  assign s_810 = s_811 & s_813;
  dq #(1, 1) dq_s_811 (clk, s_811, s_812);
  assign s_812 = s_31[23];
  assign s_813 = s_814 | s_821;
  assign s_814 = s_815 | s_817;
  dq #(1, 1) dq_s_815 (clk, s_815, s_816);
  assign s_816 = s_31[22];
  dq #(1, 1) dq_s_817 (clk, s_817, s_818);
  assign s_818 = s_819 != s_820;
  assign s_819 = s_31[21:0];
  assign s_820 = 24'd0;
  dq #(1, 1) dq_s_821 (clk, s_821, s_822);
  assign s_822 = s_30[0];
  assign s_823 = s_26[23:0];
  assign s_824 = s_26[24];
  assign s_825 = {s_826,s_837};
  assign s_826 = {s_827,s_828};
  dq #(1, 6) dq_s_827 (clk, s_827, s_3);
  assign s_828 = s_829 + s_836;
  assign s_829 = s_830[7:0];
  dq #(10, 1) dq_s_830 (clk, s_830, s_831);
  assign s_831 = s_832 + s_824;
  dq #(10, 1) dq_s_832 (clk, s_832, s_833);
  dq #(10, 1) dq_s_833 (clk, s_833, s_834);
  assign s_834 = s_835 - s_73;
  dq #(10, 2) dq_s_835 (clk, s_835, s_802);
  assign s_836 = 7'd127;
  assign s_837 = s_23[22:0];
  assign s_838 = s_839 & s_841;
  assign s_839 = s_829 == s_840;
  assign s_840 = -8'd126;
  assign s_841 = ~s_842;
  assign s_842 = s_23[23];
  assign s_843 = s_23 == s_844;
  assign s_844 = 24'd0;
  assign s_845 = s_846 | s_855;
  assign s_846 = s_847 | s_849;
  assign s_847 = $signed(s_830) > $signed(s_848);
  assign s_848 = 9'd127;
  dq #(1, 6) dq_s_849 (clk, s_849, s_850);
  assign s_850 = s_851 & s_853;
  assign s_851 = s_43 == s_852;
  assign s_852 = 8'd128;
  assign s_853 = s_47 == s_854;
  assign s_854 = 23'd0;
  dq #(1, 6) dq_s_855 (clk, s_855, s_856);
  assign s_856 = s_857 & s_859;
  assign s_857 = s_54 == s_858;
  assign s_858 = 8'd128;
  assign s_859 = s_58 == s_860;
  assign s_860 = 23'd0;
  dq #(1, 6) dq_s_861 (clk, s_861, s_862);
  assign s_862 = s_863 | s_868;
  assign s_863 = s_864 & s_866;
  assign s_864 = s_43 == s_865;
  assign s_865 = 8'd128;
  assign s_866 = s_47 != s_867;
  assign s_867 = 23'd0;
  assign s_868 = s_869 & s_871;
  assign s_869 = s_54 == s_870;
  assign s_870 = 8'd128;
  assign s_871 = s_58 != s_872;
  assign s_872 = 23'd0;
  assign mul_z = s_0;
endmodule
