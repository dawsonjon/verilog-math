//name : main_0
//input : input_data_out_1:16
//input : input_data_out_2:16
//output : output_address_1:16
//output : output_we_1:16
//output : output_data_in_1:16
//output : output_address_2:16
//output : output_we_2:16
//output : output_data_in_2:16
//source_file : fifo_tb.c

///+============================================================================+
///|                                                                            |
///|                     This file was generated by Chips                       |
///|                                                                            |
///|                                  Chips                                     |
///|                                                                            |
///|                      http://github.com/dawsonjon/Chips-2.0                 |
///|                                                                            |
///|                                                             Python powered |
///+============================================================================+
module main_0(input_data_out_1,input_data_out_2,input_data_out_1_stb,input_data_out_2_stb,output_address_1_ack,output_we_1_ack,output_data_in_1_ack,output_address_2_ack,output_we_2_ack,output_data_in_2_ack,clk,rst,output_address_1,output_we_1,output_data_in_1,output_address_2,output_we_2,output_data_in_2,output_address_1_stb,output_we_1_stb,output_data_in_1_stb,output_address_2_stb,output_we_2_stb,output_data_in_2_stb,input_data_out_1_ack,input_data_out_2_ack,exception);
  integer file_count;
  parameter  stop = 3'd0,
  instruction_fetch = 3'd1,
  operand_fetch = 3'd2,
  execute = 3'd3,
  load = 3'd4,
  wait_state = 3'd5,
  read = 3'd6,
  write = 3'd7;
  input [31:0] input_data_out_1;
  input [31:0] input_data_out_2;
  input input_data_out_1_stb;
  input input_data_out_2_stb;
  input output_address_1_ack;
  input output_we_1_ack;
  input output_data_in_1_ack;
  input output_address_2_ack;
  input output_we_2_ack;
  input output_data_in_2_ack;
  input clk;
  input rst;
  output [31:0] output_address_1;
  output [31:0] output_we_1;
  output [31:0] output_data_in_1;
  output [31:0] output_address_2;
  output [31:0] output_we_2;
  output [31:0] output_data_in_2;
  output output_address_1_stb;
  output output_we_1_stb;
  output output_data_in_1_stb;
  output output_address_2_stb;
  output output_we_2_stb;
  output output_data_in_2_stb;
  output input_data_out_1_ack;
  output input_data_out_2_ack;
  reg [31:0] timer;
  reg [63:0] timer_clock;
  reg [15:0] program_counter;
  reg [15:0] program_counter_1;
  reg [15:0] program_counter_2;
  reg [44:0] instruction;
  reg [4:0] opcode_2;
  reg [3:0] a;
  reg [3:0] b;
  reg [3:0] z;
  reg write_enable;
  reg [3:0] address_a_2;
  reg [3:0] address_b_2;
  reg [3:0] address_z_2;
  reg [3:0] address_z_3;
  reg [31:0] load_data;
  reg [31:0] write_output;
  reg [31:0] write_value;
  reg [31:0] read_input;
  reg [15:0] literal_2;
  reg [31:0] a_hi;
  reg [31:0] b_hi;
  reg [31:0] a_lo;
  reg [31:0] b_lo;
  reg [63:0] long_result;
  reg [31:0] result;
  reg [15:0] address;
  reg [31:0] data_out;
  reg [31:0] data_in;
  reg [31:0] carry;
  reg [31:0] s_output_address_1_stb;
  reg [31:0] s_output_we_1_stb;
  reg [31:0] s_output_data_in_1_stb;
  reg [31:0] s_output_address_2_stb;
  reg [31:0] s_output_we_2_stb;
  reg [31:0] s_output_data_in_2_stb;
  reg [31:0] s_output_address_1;
  reg [31:0] s_output_we_1;
  reg [31:0] s_output_data_in_1;
  reg [31:0] s_output_address_2;
  reg [31:0] s_output_we_2;
  reg [31:0] s_output_data_in_2;
  reg [31:0] s_input_data_out_1_ack;
  reg [31:0] s_input_data_out_2_ack;
  reg [7:0] state;
  output reg exception;
  reg [28:0] instructions [342:0];
  reg [31:0] memory [4096:0];
  reg [31:0] registers [15:0];
  wire [31:0] operand_a;
  wire [31:0] operand_b;
  wire [31:0] register_a;
  wire [31:0] register_b;
  wire [15:0] literal;
  wire [4:0] opcode;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] address_z;
  wire [15:0] load_address;
  wire [15:0] store_address;
  wire [31:0] store_data;
  wire  store_enable;

  //////////////////////////////////////////////////////////////////////////////
  // INSTRUCTION INITIALIZATION                                                 
  //                                                                            
  // Initialise the contents of the instruction memory                          
  //
  // Intruction Set
  // ==============
  // 0 {'literal': True, 'op': 'literal'}
  // 1 {'literal': True, 'op': 'addl'}
  // 2 {'literal': False, 'op': 'store'}
  // 3 {'literal': True, 'op': 'call'}
  // 4 {'literal': False, 'op': 'stop'}
  // 5 {'literal': False, 'op': 'load'}
  // 6 {'literal': False, 'op': 'write'}
  // 7 {'literal': False, 'op': 'greater'}
  // 8 {'literal': True, 'op': 'jmp_if_false'}
  // 9 {'literal': False, 'op': 'a_lo'}
  // 10 {'literal': False, 'line': 23, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'op': 'report'}
  // 11 {'literal': False, 'op': 'add'}
  // 12 {'literal': True, 'op': 'goto'}
  // 13 {'literal': False, 'line': 27, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'op': 'report'}
  // 14 {'literal': False, 'op': 'read'}
  // 15 {'literal': False, 'op': 'equal'}
  // 16 {'literal': False, 'line': 29, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'op': 'assert'}
  // 17 {'literal': False, 'op': 'not'}
  // 18 {'literal': False, 'line': 37, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'op': 'report'}
  // 19 {'literal': False, 'line': 41, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'op': 'report'}
  // 20 {'literal': False, 'line': 43, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'op': 'assert'}
  // 21 {'literal': False, 'op': 'return'}
  // Intructions
  // ===========
  
  initial
  begin
    instructions[0] = {5'd0, 4'd3, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46 {'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46, 'op': 'literal'}
    instructions[1] = {5'd0, 4'd4, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46 {'literal': 0, 'z': 4, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46, 'op': 'literal'}
    instructions[2] = {5'd1, 4'd3, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46 {'a': 3, 'literal': 8, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46, 'op': 'addl'}
    instructions[3] = {5'd0, 4'd8, 4'd0, 16'd2};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 3 {'literal': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 3, 'op': 'literal'}
    instructions[4] = {5'd0, 4'd2, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 3 {'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 3, 'op': 'literal'}
    instructions[5] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 3 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 3, 'op': 'store'}
    instructions[6] = {5'd0, 4'd8, 4'd0, 16'd6};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 8 {'literal': 6, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 8, 'op': 'literal'}
    instructions[7] = {5'd0, 4'd2, 4'd0, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 8 {'literal': 1, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 8, 'op': 'literal'}
    instructions[8] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 8 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 8, 'op': 'store'}
    instructions[9] = {5'd0, 4'd8, 4'd0, 16'd5};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 7 {'literal': 5, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 7, 'op': 'literal'}
    instructions[10] = {5'd0, 4'd2, 4'd0, 16'd2};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 7 {'literal': 2, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 7, 'op': 'literal'}
    instructions[11] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 7 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 7, 'op': 'store'}
    instructions[12] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 2 {'literal': 1, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 2, 'op': 'literal'}
    instructions[13] = {5'd0, 4'd2, 4'd0, 16'd3};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 2 {'literal': 3, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 2, 'op': 'literal'}
    instructions[14] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 2 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 2, 'op': 'store'}
    instructions[15] = {5'd0, 4'd8, 4'd0, 16'd4};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 6 {'literal': 4, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 6, 'op': 'literal'}
    instructions[16] = {5'd0, 4'd2, 4'd0, 16'd4};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 6 {'literal': 4, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 6, 'op': 'literal'}
    instructions[17] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 6 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 6, 'op': 'store'}
    instructions[18] = {5'd0, 4'd8, 4'd0, 16'd7};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 9 {'literal': 7, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 9, 'op': 'literal'}
    instructions[19] = {5'd0, 4'd2, 4'd0, 16'd5};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 9 {'literal': 5, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 9, 'op': 'literal'}
    instructions[20] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 9 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 9, 'op': 'store'}
    instructions[21] = {5'd0, 4'd8, 4'd0, 16'd3};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 4 {'literal': 3, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 4, 'op': 'literal'}
    instructions[22] = {5'd0, 4'd2, 4'd0, 16'd6};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 4 {'literal': 6, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 4, 'op': 'literal'}
    instructions[23] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 4 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 4, 'op': 'store'}
    instructions[24] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 1 {'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 1, 'op': 'literal'}
    instructions[25] = {5'd0, 4'd2, 4'd0, 16'd7};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 1 {'literal': 7, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 1, 'op': 'literal'}
    instructions[26] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 1 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 1, 'op': 'store'}
    instructions[27] = {5'd1, 4'd7, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46 {'a': 4, 'literal': 0, 'z': 7, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46, 'op': 'addl'}
    instructions[28] = {5'd1, 4'd4, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46 {'a': 3, 'literal': 0, 'z': 4, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46, 'op': 'addl'}
    instructions[29] = {5'd3, 4'd6, 4'd0, 16'd31};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46 {'z': 6, 'label': 31, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46, 'op': 'call'}
    instructions[30] = {5'd4, 4'd0, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46 {'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 46, 'op': 'stop'}
    instructions[31] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 11 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 11, 'op': 'addl'}
    instructions[32] = {5'd0, 4'd8, 4'd0, 16'd3};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14 {'literal': 3, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14, 'op': 'literal'}
    instructions[33] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14, 'op': 'addl'}
    instructions[34] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14, 'op': 'load'}
    instructions[35] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14, 'op': 'store'}
    instructions[36] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14, 'op': 'addl'}
    instructions[37] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14 {'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14, 'op': 'literal'}
    instructions[38] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[39] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14, 'op': 'load'}
    instructions[40] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14, 'op': 'write'}
    instructions[41] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 14, 'op': 'addl'}
    instructions[42] = {5'd0, 4'd8, 4'd0, 16'd2};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15 {'literal': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15, 'op': 'literal'}
    instructions[43] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15, 'op': 'addl'}
    instructions[44] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15, 'op': 'load'}
    instructions[45] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15, 'op': 'store'}
    instructions[46] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15, 'op': 'addl'}
    instructions[47] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15 {'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15, 'op': 'literal'}
    instructions[48] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[49] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15, 'op': 'load'}
    instructions[50] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15, 'op': 'write'}
    instructions[51] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 15, 'op': 'addl'}
    instructions[52] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'literal'}
    instructions[53] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[54] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'store'}
    instructions[55] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[56] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[57] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'load'}
    instructions[58] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'store'}
    instructions[59] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[60] = {5'd0, 4'd8, 4'd0, 16'd256};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'literal': 256, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'literal'}
    instructions[61] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[62] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'z': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'load'}
    instructions[63] = {5'd7, 4'd8, 4'd8, 16'd10};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'greater'}
    instructions[64] = {5'd8, 4'd0, 4'd8, 16'd133};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 8, 'label': 133, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'jmp_if_false'}
    instructions[65] = {5'd0, 4'd8, 4'd0, 16'd7};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'literal': 7, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'literal'}
    instructions[66] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'addl'}
    instructions[67] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'load'}
    instructions[68] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'store'}
    instructions[69] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'addl'}
    instructions[70] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'addl'}
    instructions[71] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'addl'}
    instructions[72] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'load'}
    instructions[73] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[74] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'load'}
    instructions[75] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'write'}
    instructions[76] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 18, 'op': 'addl'}
    instructions[77] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'literal'}
    instructions[78] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'addl'}
    instructions[79] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'load'}
    instructions[80] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'store'}
    instructions[81] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'addl'}
    instructions[82] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'addl'}
    instructions[83] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'addl'}
    instructions[84] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'load'}
    instructions[85] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[86] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'load'}
    instructions[87] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'write'}
    instructions[88] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 19, 'op': 'addl'}
    instructions[89] = {5'd0, 4'd8, 4'd0, 16'd3};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20 {'literal': 3, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20, 'op': 'literal'}
    instructions[90] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20, 'op': 'addl'}
    instructions[91] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20, 'op': 'load'}
    instructions[92] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20, 'op': 'store'}
    instructions[93] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20, 'op': 'addl'}
    instructions[94] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20 {'literal': 1, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20, 'op': 'literal'}
    instructions[95] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[96] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20, 'op': 'load'}
    instructions[97] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20, 'op': 'write'}
    instructions[98] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 20, 'op': 'addl'}
    instructions[99] = {5'd0, 4'd8, 4'd0, 16'd3};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21 {'literal': 3, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21, 'op': 'literal'}
    instructions[100] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21, 'op': 'addl'}
    instructions[101] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21, 'op': 'load'}
    instructions[102] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21, 'op': 'store'}
    instructions[103] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21, 'op': 'addl'}
    instructions[104] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21 {'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21, 'op': 'literal'}
    instructions[105] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[106] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21, 'op': 'load'}
    instructions[107] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21, 'op': 'write'}
    instructions[108] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 21, 'op': 'addl'}
    instructions[109] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 22 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 22, 'op': 'addl'}
    instructions[110] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 22 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 22, 'op': 'addl'}
    instructions[111] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 22 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 22, 'op': 'load'}
    instructions[112] = {5'd9, 4'd8, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 22 {'a': 8, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 22, 'op': 'a_lo'}
    instructions[113] = {5'd10, 4'd0, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 22 {'line': 23, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 22, 'op': 'report'}
    instructions[114] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[115] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[116] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'load'}
    instructions[117] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'store'}
    instructions[118] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[119] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'literal': 1, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'literal'}
    instructions[120] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'store'}
    instructions[121] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[122] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[123] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[124] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'load'}
    instructions[125] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[126] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'z': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'load'}
    instructions[127] = {5'd11, 4'd8, 4'd8, 16'd10};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'add'}
    instructions[128] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'addl'}
    instructions[129] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'store'}
    instructions[130] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[131] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'a': 3, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'load'}
    instructions[132] = {5'd12, 4'd0, 4'd0, 16'd55};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17 {'label': 55, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 17, 'op': 'goto'}
    instructions[133] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'literal'}
    instructions[134] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[135] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'store'}
    instructions[136] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[137] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[138] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'load'}
    instructions[139] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'store'}
    instructions[140] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[141] = {5'd0, 4'd8, 4'd0, 16'd256};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'literal': 256, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'literal'}
    instructions[142] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[143] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'z': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'load'}
    instructions[144] = {5'd7, 4'd8, 4'd8, 16'd10};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'greater'}
    instructions[145] = {5'd8, 4'd0, 4'd8, 16'd195};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 8, 'label': 195, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'jmp_if_false'}
    instructions[146] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 26 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 26, 'op': 'addl'}
    instructions[147] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 26 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 26, 'op': 'addl'}
    instructions[148] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 26 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 26, 'op': 'load'}
    instructions[149] = {5'd9, 4'd8, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 26 {'a': 8, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 26, 'op': 'a_lo'}
    instructions[150] = {5'd13, 4'd0, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 26 {'line': 27, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 26, 'op': 'report'}
    instructions[151] = {5'd0, 4'd8, 4'd0, 16'd4};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'literal': 4, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'literal'}
    instructions[152] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'addl'}
    instructions[153] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'load'}
    instructions[154] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'store'}
    instructions[155] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'addl'}
    instructions[156] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'addl'}
    instructions[157] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'addl'}
    instructions[158] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'load'}
    instructions[159] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[160] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'load'}
    instructions[161] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'write'}
    instructions[162] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 27, 'op': 'addl'}
    instructions[163] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'addl'}
    instructions[164] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'addl'}
    instructions[165] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'load'}
    instructions[166] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'store'}
    instructions[167] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'addl'}
    instructions[168] = {5'd0, 4'd8, 4'd0, 16'd5};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'literal': 5, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'literal'}
    instructions[169] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'addl'}
    instructions[170] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'load'}
    instructions[171] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 8, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'read'}
    instructions[172] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[173] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 3, 'z': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'load'}
    instructions[174] = {5'd15, 4'd8, 4'd8, 16'd10};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'equal'}
    instructions[175] = {5'd16, 4'd0, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28 {'a': 8, 'line': 29, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 28, 'op': 'assert'}
    instructions[176] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[177] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[178] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'load'}
    instructions[179] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'store'}
    instructions[180] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[181] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'literal': 1, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'literal'}
    instructions[182] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'store'}
    instructions[183] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[184] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[185] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[186] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'load'}
    instructions[187] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[188] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'z': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'load'}
    instructions[189] = {5'd11, 4'd8, 4'd8, 16'd10};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'add'}
    instructions[190] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'addl'}
    instructions[191] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'store'}
    instructions[192] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[193] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'a': 3, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'load'}
    instructions[194] = {5'd12, 4'd0, 4'd0, 16'd136};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25 {'label': 136, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 25, 'op': 'goto'}
    instructions[195] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'literal'}
    instructions[196] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[197] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'store'}
    instructions[198] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[199] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[200] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'load'}
    instructions[201] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'store'}
    instructions[202] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[203] = {5'd0, 4'd8, 4'd0, 16'd256};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'literal': 256, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'literal'}
    instructions[204] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[205] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'z': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'load'}
    instructions[206] = {5'd7, 4'd8, 4'd8, 16'd10};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'greater'}
    instructions[207] = {5'd8, 4'd0, 4'd8, 16'd277};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 8, 'label': 277, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'jmp_if_false'}
    instructions[208] = {5'd0, 4'd8, 4'd0, 16'd4};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'literal': 4, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'literal'}
    instructions[209] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'addl'}
    instructions[210] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'load'}
    instructions[211] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'store'}
    instructions[212] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'addl'}
    instructions[213] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'addl'}
    instructions[214] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'addl'}
    instructions[215] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'load'}
    instructions[216] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[217] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'load'}
    instructions[218] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'write'}
    instructions[219] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 32, 'op': 'addl'}
    instructions[220] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'literal': 1, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'literal'}
    instructions[221] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'addl'}
    instructions[222] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'load'}
    instructions[223] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'store'}
    instructions[224] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'addl'}
    instructions[225] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'addl'}
    instructions[226] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'addl'}
    instructions[227] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'load'}
    instructions[228] = {5'd17, 4'd8, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 8, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'not'}
    instructions[229] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[230] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'load'}
    instructions[231] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'write'}
    instructions[232] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 33, 'op': 'addl'}
    instructions[233] = {5'd0, 4'd8, 4'd0, 16'd2};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34 {'literal': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34, 'op': 'literal'}
    instructions[234] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34, 'op': 'addl'}
    instructions[235] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34, 'op': 'load'}
    instructions[236] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34, 'op': 'store'}
    instructions[237] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34, 'op': 'addl'}
    instructions[238] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34 {'literal': 1, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34, 'op': 'literal'}
    instructions[239] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[240] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34, 'op': 'load'}
    instructions[241] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34, 'op': 'write'}
    instructions[242] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 34, 'op': 'addl'}
    instructions[243] = {5'd0, 4'd8, 4'd0, 16'd2};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35 {'literal': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35, 'op': 'literal'}
    instructions[244] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35, 'op': 'addl'}
    instructions[245] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35, 'op': 'load'}
    instructions[246] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35, 'op': 'store'}
    instructions[247] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35, 'op': 'addl'}
    instructions[248] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35 {'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35, 'op': 'literal'}
    instructions[249] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[250] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35, 'op': 'load'}
    instructions[251] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35, 'op': 'write'}
    instructions[252] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 35, 'op': 'addl'}
    instructions[253] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 36 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 36, 'op': 'addl'}
    instructions[254] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 36 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 36, 'op': 'addl'}
    instructions[255] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 36 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 36, 'op': 'load'}
    instructions[256] = {5'd9, 4'd8, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 36 {'a': 8, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 36, 'op': 'a_lo'}
    instructions[257] = {5'd18, 4'd0, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 36 {'line': 37, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 36, 'op': 'report'}
    instructions[258] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[259] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[260] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'load'}
    instructions[261] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'store'}
    instructions[262] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[263] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'literal': 1, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'literal'}
    instructions[264] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'store'}
    instructions[265] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[266] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[267] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[268] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'load'}
    instructions[269] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[270] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'z': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'load'}
    instructions[271] = {5'd11, 4'd8, 4'd8, 16'd10};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'add'}
    instructions[272] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'addl'}
    instructions[273] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'store'}
    instructions[274] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[275] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'a': 3, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'load'}
    instructions[276] = {5'd12, 4'd0, 4'd0, 16'd198};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31 {'label': 198, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 31, 'op': 'goto'}
    instructions[277] = {5'd0, 4'd8, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'literal'}
    instructions[278] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[279] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'store'}
    instructions[280] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[281] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[282] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'load'}
    instructions[283] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'store'}
    instructions[284] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[285] = {5'd0, 4'd8, 4'd0, 16'd256};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'literal': 256, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'literal'}
    instructions[286] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[287] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'z': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'load'}
    instructions[288] = {5'd7, 4'd8, 4'd8, 16'd10};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'greater'}
    instructions[289] = {5'd8, 4'd0, 4'd8, 16'd340};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 8, 'label': 340, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'jmp_if_false'}
    instructions[290] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 40 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 40, 'op': 'addl'}
    instructions[291] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 40 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 40, 'op': 'addl'}
    instructions[292] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 40 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 40, 'op': 'load'}
    instructions[293] = {5'd9, 4'd8, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 40 {'a': 8, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 40, 'op': 'a_lo'}
    instructions[294] = {5'd19, 4'd0, 4'd0, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 40 {'line': 41, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 40, 'op': 'report'}
    instructions[295] = {5'd0, 4'd8, 4'd0, 16'd7};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'literal': 7, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'literal'}
    instructions[296] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'addl'}
    instructions[297] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'load'}
    instructions[298] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'store'}
    instructions[299] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'addl'}
    instructions[300] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'addl'}
    instructions[301] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'addl'}
    instructions[302] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'load'}
    instructions[303] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[304] = {5'd5, 4'd0, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 3, 'z': 0, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'load'}
    instructions[305] = {5'd6, 4'd0, 4'd0, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 0, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'write'}
    instructions[306] = {5'd1, 4'd3, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41 {'a': 3, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 41, 'op': 'addl'}
    instructions[307] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'addl'}
    instructions[308] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'addl'}
    instructions[309] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'load'}
    instructions[310] = {5'd17, 4'd8, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 8, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'not'}
    instructions[311] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'store'}
    instructions[312] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'addl'}
    instructions[313] = {5'd0, 4'd8, 4'd0, 16'd6};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'literal': 6, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'literal'}
    instructions[314] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'addl'}
    instructions[315] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'load'}
    instructions[316] = {5'd14, 4'd8, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 8, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'read'}
    instructions[317] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[318] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 3, 'z': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'load'}
    instructions[319] = {5'd15, 4'd8, 4'd8, 16'd10};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'equal'}
    instructions[320] = {5'd20, 4'd0, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42 {'a': 8, 'line': 43, 'file': '/home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 42, 'op': 'assert'}
    instructions[321] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[322] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[323] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'load'}
    instructions[324] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'store'}
    instructions[325] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[326] = {5'd0, 4'd8, 4'd0, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'literal': 1, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'literal'}
    instructions[327] = {5'd2, 4'd0, 4'd3, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'comment': 'push', 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'store'}
    instructions[328] = {5'd1, 4'd3, 4'd3, 16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'literal': 1, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[329] = {5'd1, 4'd8, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 4, 'literal': 0, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[330] = {5'd1, 4'd2, 4'd8, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 8, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[331] = {5'd5, 4'd8, 4'd2, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 2, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'load'}
    instructions[332] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[333] = {5'd5, 4'd10, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'z': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'load'}
    instructions[334] = {5'd11, 4'd8, 4'd8, 16'd10};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 8, 'z': 8, 'b': 10, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'add'}
    instructions[335] = {5'd1, 4'd2, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 4, 'literal': 0, 'z': 2, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'addl'}
    instructions[336] = {5'd2, 4'd0, 4'd2, 16'd8};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 2, 'b': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'store'}
    instructions[337] = {5'd1, 4'd3, 4'd3, -16'd1};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'comment': 'pop', 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'literal': -1, 'z': 3, 'op': 'addl'}
    instructions[338] = {5'd5, 4'd8, 4'd3, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'a': 3, 'z': 8, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'load'}
    instructions[339] = {5'd12, 4'd0, 4'd0, 16'd280};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39 {'label': 280, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 39, 'op': 'goto'}
    instructions[340] = {5'd1, 4'd3, 4'd4, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 11 {'a': 4, 'literal': 0, 'z': 3, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 11, 'op': 'addl'}
    instructions[341] = {5'd1, 4'd4, 4'd7, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 11 {'a': 7, 'literal': 0, 'z': 4, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 11, 'op': 'addl'}
    instructions[342] = {5'd21, 4'd0, 4'd6, 16'd0};///home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 11 {'a': 6, 'trace': /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c : 11, 'op': 'return'}
  end

  
  always @(posedge clk)
  begin
    load_data <= memory[load_address];
    if(store_enable && state == execute) begin
      memory[store_address] <= store_data;
    end
  end


  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 1 -- FETCH INSTRUCTION
  //                                                                            
  
  always @(posedge clk)
  begin
    //implement memory for instructions
    if (state == instruction_fetch || state == operand_fetch || state == execute) begin
      instruction <= instructions[program_counter];
      program_counter_1 <= program_counter;
    end
  end

  assign opcode    = instruction[28:24];
  assign address_z = instruction[23:20];
  assign address_a = instruction[19:16];
  assign address_b = instruction[3:0];
  assign literal   = instruction[15:0];

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 2 -- FETCH OPERANDS
  //                                                                            
  
  always @(posedge clk)
  begin
    if (write_enable) begin
      registers[address_z_3] <= result;
    end
    if (state == operand_fetch || state == execute) begin
      opcode_2 <= opcode;
      literal_2 <= literal;
      address_a_2 <= address_a;
      address_b_2 <= address_b;
      address_z_2 <= address_z;
      program_counter_2 <= program_counter_1;
    end
  end
  assign register_a = registers[address_a_2];
  assign register_b = registers[address_b_2];
  assign operand_a = (address_a_2 == address_z_3 && write_enable)?result:register_a;
  assign operand_b = (address_b_2 == address_z_3 && write_enable)?result:register_b;
  assign store_address = operand_a;
  assign load_address = operand_a;
  assign store_data = operand_b;
  assign store_enable = (opcode_2==2);

  //////////////////////////////////////////////////////////////////////////////
  // PIPELINE STAGE 3 -- EXECUTE
  //                                                                            
  
  always @(posedge clk)
  begin

  write_enable <= 0;
  timer_clock <= timer_clock + 1;
  case(state)

    //instruction_fetch
    instruction_fetch: begin
      program_counter <= program_counter + 1;
      state <= operand_fetch;
    end
    //operand_fetch
    operand_fetch: begin
      program_counter <= program_counter + 1;
      state <= execute;
    end
    //execute
    execute: begin
      program_counter <= program_counter + 1;
      address_z_3 <= address_z_2;
      case(opcode_2)

        //literal
        16'd0:
        begin
          result<=$signed(literal_2);
          write_enable <= 1;
        end

        //addl
        16'd1:
        begin
          result<=operand_a + literal_2;
          write_enable <= 1;
        end

        //store
        16'd2:
        begin
        end

        //call
        16'd3:
        begin
          result <= program_counter_2 + 1;
          write_enable <= 1;
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //stop
        16'd4:
        begin
        state <= stop;
        end

        //load
        16'd5:
        begin
          state <= load;
        end

        //write
        16'd6:
        begin
          state <= write;
          write_output <= operand_a;
          write_value <= operand_b;
        end

        //greater
        16'd7:
        begin
          result <= $signed(operand_a) > $signed(operand_b);
          write_enable <= 1;
        end

        //jmp_if_false
        16'd8:
        begin
          if (operand_a == 0) begin
            program_counter <= literal_2;
            state <= instruction_fetch;
          end
        end

        //a_lo
        16'd9:
        begin
          a_lo <= operand_a;
          result <= a_lo;
          write_enable <= 1;
        end

        //report
        16'd10:
        begin
          $display ("%d (report (int) at line: 23 in file: /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c)", $signed(a_lo));
        end

        //add
        16'd11:
        begin
          long_result = operand_a + operand_b;
          result <= long_result[31:0];
          carry[0] <= long_result[32];
          write_enable <= 1;
        end

        //goto
        16'd12:
        begin
          program_counter <= literal_2;
          state <= instruction_fetch;
        end

        //report
        16'd13:
        begin
          $display ("%d (report (int) at line: 27 in file: /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c)", $signed(a_lo));
        end

        //read
        16'd14:
        begin
          state <= read;
          read_input <= operand_a;
        end

        //equal
        16'd15:
        begin
          result <= operand_a == operand_b;
          write_enable <= 1;
        end

        //assert
        16'd16:
        begin
          if (operand_a == 0) begin
            $display("Assertion failed at line: 29 in file: /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c");
            $finish_and_return(1);
          end
        end

        //not
        16'd17:
        begin
          result <= ~operand_a;
          write_enable <= 1;
        end

        //report
        16'd18:
        begin
          $display ("%d (report (int) at line: 37 in file: /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c)", $signed(a_lo));
        end

        //report
        16'd19:
        begin
          $display ("%d (report (int) at line: 41 in file: /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c)", $signed(a_lo));
        end

        //assert
        16'd20:
        begin
          if (operand_a == 0) begin
            $display("Assertion failed at line: 43 in file: /home/jon/portable_ip_library/components/memory/fifo/test/fifo_tb.c");
            $finish_and_return(1);
          end
        end

        //return
        16'd21:
        begin
          program_counter <= operand_a;
          state <= instruction_fetch;
        end

      endcase

    end

    read:
    begin
      case(read_input)
      3:
      begin
        s_input_data_out_1_ack <= 1;
        if (s_input_data_out_1_ack && input_data_out_1_stb) begin
          result <= input_data_out_1;
          write_enable <= 1;
          s_input_data_out_1_ack <= 0;
          state <= execute;
        end
      end
      7:
      begin
        s_input_data_out_2_ack <= 1;
        if (s_input_data_out_2_ack && input_data_out_2_stb) begin
          result <= input_data_out_2;
          write_enable <= 1;
          s_input_data_out_2_ack <= 0;
          state <= execute;
        end
      end
      endcase
    end

    write:
    begin
      case(write_output)
      0:
      begin
        s_output_address_1_stb <= 1;
        s_output_address_1 <= write_value;
        if (output_address_1_ack && s_output_address_1_stb) begin
          s_output_address_1_stb <= 0;
          state <= execute;
        end
      end
      1:
      begin
        s_output_we_1_stb <= 1;
        s_output_we_1 <= write_value;
        if (output_we_1_ack && s_output_we_1_stb) begin
          s_output_we_1_stb <= 0;
          state <= execute;
        end
      end
      2:
      begin
        s_output_data_in_1_stb <= 1;
        s_output_data_in_1 <= write_value;
        if (output_data_in_1_ack && s_output_data_in_1_stb) begin
          s_output_data_in_1_stb <= 0;
          state <= execute;
        end
      end
      4:
      begin
        s_output_address_2_stb <= 1;
        s_output_address_2 <= write_value;
        if (output_address_2_ack && s_output_address_2_stb) begin
          s_output_address_2_stb <= 0;
          state <= execute;
        end
      end
      5:
      begin
        s_output_we_2_stb <= 1;
        s_output_we_2 <= write_value;
        if (output_we_2_ack && s_output_we_2_stb) begin
          s_output_we_2_stb <= 0;
          state <= execute;
        end
      end
      6:
      begin
        s_output_data_in_2_stb <= 1;
        s_output_data_in_2 <= write_value;
        if (output_data_in_2_ack && s_output_data_in_2_stb) begin
          s_output_data_in_2_stb <= 0;
          state <= execute;
        end
      end
      endcase
    end

    load:
    begin
        result <= load_data;
        write_enable <= 1;
        state <= execute;
    end

    wait_state:
    begin
      if (timer) begin
        timer <= timer - 1;
      end else begin
        state <= execute;
      end
    end

    stop:
    begin
    end

    endcase

    if (rst == 1'b1) begin
      timer <= 0;
      timer_clock <= 0;
      program_counter <= 0;
      address_z_3 <= 0;
      result <= 0;
      a = 0;
      b = 0;
      z = 0;
      state <= instruction_fetch;
      s_input_data_out_1_ack <= 0;
      s_input_data_out_2_ack <= 0;
      s_output_address_1_stb <= 0;
      s_output_we_1_stb <= 0;
      s_output_data_in_1_stb <= 0;
      s_output_address_2_stb <= 0;
      s_output_we_2_stb <= 0;
      s_output_data_in_2_stb <= 0;
    end
  end
  assign input_data_out_1_ack = s_input_data_out_1_ack;
  assign input_data_out_2_ack = s_input_data_out_2_ack;
  assign output_address_1_stb = s_output_address_1_stb;
  assign output_address_1 = s_output_address_1;
  assign output_we_1_stb = s_output_we_1_stb;
  assign output_we_1 = s_output_we_1;
  assign output_data_in_1_stb = s_output_data_in_1_stb;
  assign output_data_in_1 = s_output_data_in_1;
  assign output_address_2_stb = s_output_address_2_stb;
  assign output_address_2 = s_output_address_2;
  assign output_we_2_stb = s_output_we_2_stb;
  assign output_we_2 = s_output_we_2;
  assign output_data_in_2_stb = s_output_data_in_2_stb;
  assign output_data_in_2 = s_output_data_in_2;

endmodule
