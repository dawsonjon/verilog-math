module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module ne(clk, ne_a, ne_b, ne_z);
  input clk;
  input [31:0] ne_a;
  input [31:0] ne_b;
  output [0:0] ne_z;
  wire [0:0] s_0;
  wire [0:0] s_1;
  wire [0:0] s_2;
  wire [0:0] s_3;
  wire [0:0] s_4;
  wire [0:0] s_5;
  wire [31:0] s_6;
  wire [0:0] s_7;
  wire [31:0] s_8;
  wire [0:0] s_9;
  wire [7:0] s_10;
  wire [7:0] s_11;
  wire [7:0] s_12;
  wire [7:0] s_13;
  wire [6:0] s_14;
  wire [0:0] s_15;
  wire [7:0] s_16;
  wire [7:0] s_17;
  wire [7:0] s_18;
  wire [7:0] s_19;
  wire [7:0] s_20;
  wire [6:0] s_21;
  wire [0:0] s_22;
  wire [7:0] s_23;
  wire [0:0] s_24;
  wire [23:0] s_25;
  wire [0:0] s_26;
  wire [0:0] s_27;
  wire [0:0] s_28;
  wire [22:0] s_29;
  wire [23:0] s_30;
  wire [0:0] s_31;
  wire [0:0] s_32;
  wire [0:0] s_33;
  wire [22:0] s_34;
  wire [0:0] s_35;
  wire [0:0] s_36;
  wire [0:0] s_37;
  wire [0:0] s_38;
  wire [0:0] s_39;
  wire [0:0] s_40;
  wire [0:0] s_41;
  wire [0:0] s_42;
  wire [0:0] s_43;
  wire [0:0] s_44;
  wire [0:0] s_45;
  wire [7:0] s_46;
  wire [0:0] s_47;
  wire [22:0] s_48;
  wire [0:0] s_49;
  wire [0:0] s_50;
  wire [0:0] s_51;
  wire [7:0] s_52;
  wire [0:0] s_53;
  wire [22:0] s_54;

  assign s_0 = ~s_1;
  assign s_1 = s_2 | s_35;
  assign s_2 = s_3 & s_24;
  assign s_3 = s_4 & s_9;
  assign s_4 = s_5 == s_7;
  assign s_5 = s_6[31];
  assign s_6 = ne_a;
  assign s_7 = s_8[31];
  assign s_8 = ne_b;
  assign s_9 = s_10 == s_17;
  assign s_10 = s_15?s_11:s_12;
  assign s_11 = -8'd126;
  assign s_12 = s_13 - s_14;
  assign s_13 = s_6[30:23];
  assign s_14 = 7'd127;
  assign s_15 = s_12 == s_16;
  assign s_16 = -8'd127;
  assign s_17 = s_22?s_18:s_19;
  assign s_18 = -8'd126;
  assign s_19 = s_20 - s_21;
  assign s_20 = s_8[30:23];
  assign s_21 = 7'd127;
  assign s_22 = s_19 == s_23;
  assign s_23 = -8'd127;
  assign s_24 = s_25 == s_30;
  assign s_25 = {s_26,s_29};
  assign s_26 = s_15?s_27:s_28;
  assign s_27 = 1'd0;
  assign s_28 = 1'd1;
  assign s_29 = s_6[22:0];
  assign s_30 = {s_31,s_34};
  assign s_31 = s_22?s_32:s_33;
  assign s_32 = 1'd0;
  assign s_33 = 1'd1;
  assign s_34 = s_8[22:0];
  assign s_35 = s_36 & s_49;
  assign s_36 = s_37 & s_43;
  assign s_37 = s_38 & s_41;
  assign s_38 = s_39 & s_40;
  assign s_39 = s_10 == s_17;
  assign s_40 = s_25 == s_30;
  assign s_41 = s_25 == s_42;
  assign s_42 = 1'd0;
  assign s_43 = ~s_44;
  assign s_44 = s_45 & s_47;
  assign s_45 = s_12 == s_46;
  assign s_46 = 8'd128;
  assign s_47 = s_29 != s_48;
  assign s_48 = 23'd0;
  assign s_49 = ~s_50;
  assign s_50 = s_51 & s_53;
  assign s_51 = s_19 == s_52;
  assign s_52 = 8'd128;
  assign s_53 = s_34 != s_54;
  assign s_54 = 23'd0;
  assign ne_z = s_0;
endmodule
