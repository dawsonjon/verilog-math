module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module double_add(clk, double_add_a, double_add_b, double_add_z);
  input clk;
  input [63:0] double_add_a;
  input [63:0] double_add_b;
  output [63:0] double_add_z;
  wire [63:0] s_0;
  wire [63:0] s_1;
  wire [63:0] s_2;
  wire [0:0] s_3;
  wire [0:0] s_4;
  wire [0:0] s_5;
  wire [0:0] s_6;
  wire [0:0] s_7;
  wire [0:0] s_8;
  wire [63:0] s_9;
  wire [0:0] s_10;
  wire [63:0] s_11;
  wire [0:0] s_12;
  wire [0:0] s_13;
  wire [0:0] s_14;
  wire [11:0] s_15;
  wire [10:0] s_16;
  wire [10:0] s_17;
  wire [10:0] s_18;
  wire [10:0] s_19;
  wire [9:0] s_20;
  wire [0:0] s_21;
  wire [10:0] s_22;
  wire [11:0] s_23;
  wire [10:0] s_24;
  wire [10:0] s_25;
  wire [10:0] s_26;
  wire [10:0] s_27;
  wire [9:0] s_28;
  wire [0:0] s_29;
  wire [10:0] s_30;
  wire [0:0] s_31;
  wire [0:0] s_32;
  wire [10:0] s_33;
  wire [0:0] s_34;
  wire [51:0] s_35;
  wire [51:0] s_36;
  wire [0:0] s_37;
  wire [0:0] s_38;
  wire [0:0] s_39;
  wire [10:0] s_40;
  wire [0:0] s_41;
  wire [51:0] s_42;
  wire [51:0] s_43;
  wire [0:0] s_44;
  wire [0:0] s_45;
  wire [56:0] s_46;
  wire [56:0] s_47;
  wire [52:0] s_48;
  wire [52:0] s_49;
  wire [0:0] s_50;
  wire [0:0] s_51;
  wire [0:0] s_52;
  wire [52:0] s_53;
  wire [0:0] s_54;
  wire [0:0] s_55;
  wire [0:0] s_56;
  wire [1:0] s_57;
  wire [56:0] s_58;
  wire [56:0] s_59;
  wire [56:0] s_60;
  wire [56:0] s_61;
  wire [52:0] s_62;
  wire [1:0] s_63;
  wire [11:0] s_64;
  wire [11:0] s_65;
  wire [11:0] s_66;
  wire [0:0] s_67;
  wire [56:0] s_68;
  wire [56:0] s_69;
  wire [56:0] s_70;
  wire [0:0] s_71;
  wire [0:0] s_72;
  wire [56:0] s_73;
  wire [56:0] s_74;
  wire [56:0] s_75;
  wire [56:0] s_76;
  wire [56:0] s_77;
  wire [56:0] s_78;
  wire [56:0] s_79;
  wire [56:0] s_80;
  wire [56:0] s_81;
  wire [0:0] s_82;
  wire [0:0] s_83;
  wire [62:0] s_84;
  wire [63:0] s_85;
  wire [63:0] s_86;
  wire [63:0] s_87;
  wire [62:0] s_88;
  wire [63:0] s_89;
  wire [63:0] s_90;
  wire [63:0] s_91;
  wire [62:0] s_92;
  wire [63:0] s_93;
  wire [63:0] s_94;
  wire [11:0] s_95;
  wire [11:0] s_96;
  wire [10:0] s_97;
  wire [51:0] s_98;
  wire [52:0] s_99;
  wire [52:0] s_100;
  wire [52:0] s_101;
  wire [53:0] s_102;
  wire [53:0] s_103;
  wire [53:0] s_104;
  wire [53:0] s_105;
  wire [52:0] s_106;
  wire [56:0] s_107;
  wire [56:0] s_108;
  wire [56:0] s_109;
  wire [56:0] s_110;
  wire [11:0] s_111;
  wire [11:0] s_112;
  wire [6:0] s_113;
  wire [6:0] s_114;
  wire [0:0] s_115;
  wire [0:0] s_116;
  wire [5:0] s_117;
  wire [0:0] s_118;
  wire [0:0] s_119;
  wire [4:0] s_120;
  wire [0:0] s_121;
  wire [0:0] s_122;
  wire [3:0] s_123;
  wire [0:0] s_124;
  wire [0:0] s_125;
  wire [2:0] s_126;
  wire [0:0] s_127;
  wire [0:0] s_128;
  wire [1:0] s_129;
  wire [0:0] s_130;
  wire [0:0] s_131;
  wire [0:0] s_132;
  wire [1:0] s_133;
  wire [3:0] s_134;
  wire [7:0] s_135;
  wire [15:0] s_136;
  wire [31:0] s_137;
  wire [63:0] s_138;
  wire [62:0] s_139;
  wire [61:0] s_140;
  wire [60:0] s_141;
  wire [59:0] s_142;
  wire [58:0] s_143;
  wire [57:0] s_144;
  wire [0:0] s_145;
  wire [0:0] s_146;
  wire [0:0] s_147;
  wire [0:0] s_148;
  wire [0:0] s_149;
  wire [0:0] s_150;
  wire [0:0] s_151;
  wire [0:0] s_152;
  wire [0:0] s_153;
  wire [0:0] s_154;
  wire [0:0] s_155;
  wire [0:0] s_156;
  wire [0:0] s_157;
  wire [0:0] s_158;
  wire [1:0] s_159;
  wire [0:0] s_160;
  wire [0:0] s_161;
  wire [0:0] s_162;
  wire [1:0] s_163;
  wire [0:0] s_164;
  wire [0:0] s_165;
  wire [0:0] s_166;
  wire [0:0] s_167;
  wire [0:0] s_168;
  wire [0:0] s_169;
  wire [1:0] s_170;
  wire [0:0] s_171;
  wire [0:0] s_172;
  wire [0:0] s_173;
  wire [0:0] s_174;
  wire [0:0] s_175;
  wire [0:0] s_176;
  wire [2:0] s_177;
  wire [0:0] s_178;
  wire [0:0] s_179;
  wire [1:0] s_180;
  wire [0:0] s_181;
  wire [0:0] s_182;
  wire [0:0] s_183;
  wire [1:0] s_184;
  wire [3:0] s_185;
  wire [0:0] s_186;
  wire [0:0] s_187;
  wire [0:0] s_188;
  wire [0:0] s_189;
  wire [0:0] s_190;
  wire [0:0] s_191;
  wire [0:0] s_192;
  wire [1:0] s_193;
  wire [0:0] s_194;
  wire [0:0] s_195;
  wire [0:0] s_196;
  wire [1:0] s_197;
  wire [0:0] s_198;
  wire [0:0] s_199;
  wire [0:0] s_200;
  wire [0:0] s_201;
  wire [0:0] s_202;
  wire [0:0] s_203;
  wire [1:0] s_204;
  wire [0:0] s_205;
  wire [0:0] s_206;
  wire [0:0] s_207;
  wire [0:0] s_208;
  wire [0:0] s_209;
  wire [2:0] s_210;
  wire [0:0] s_211;
  wire [0:0] s_212;
  wire [1:0] s_213;
  wire [1:0] s_214;
  wire [1:0] s_215;
  wire [0:0] s_216;
  wire [3:0] s_217;
  wire [0:0] s_218;
  wire [0:0] s_219;
  wire [2:0] s_220;
  wire [0:0] s_221;
  wire [0:0] s_222;
  wire [1:0] s_223;
  wire [0:0] s_224;
  wire [0:0] s_225;
  wire [0:0] s_226;
  wire [1:0] s_227;
  wire [3:0] s_228;
  wire [7:0] s_229;
  wire [0:0] s_230;
  wire [0:0] s_231;
  wire [0:0] s_232;
  wire [0:0] s_233;
  wire [0:0] s_234;
  wire [0:0] s_235;
  wire [0:0] s_236;
  wire [1:0] s_237;
  wire [0:0] s_238;
  wire [0:0] s_239;
  wire [0:0] s_240;
  wire [1:0] s_241;
  wire [0:0] s_242;
  wire [0:0] s_243;
  wire [0:0] s_244;
  wire [0:0] s_245;
  wire [0:0] s_246;
  wire [0:0] s_247;
  wire [1:0] s_248;
  wire [0:0] s_249;
  wire [0:0] s_250;
  wire [0:0] s_251;
  wire [0:0] s_252;
  wire [0:0] s_253;
  wire [0:0] s_254;
  wire [2:0] s_255;
  wire [0:0] s_256;
  wire [0:0] s_257;
  wire [1:0] s_258;
  wire [0:0] s_259;
  wire [0:0] s_260;
  wire [0:0] s_261;
  wire [1:0] s_262;
  wire [3:0] s_263;
  wire [0:0] s_264;
  wire [0:0] s_265;
  wire [0:0] s_266;
  wire [0:0] s_267;
  wire [0:0] s_268;
  wire [0:0] s_269;
  wire [0:0] s_270;
  wire [1:0] s_271;
  wire [0:0] s_272;
  wire [0:0] s_273;
  wire [0:0] s_274;
  wire [1:0] s_275;
  wire [0:0] s_276;
  wire [0:0] s_277;
  wire [0:0] s_278;
  wire [0:0] s_279;
  wire [0:0] s_280;
  wire [0:0] s_281;
  wire [1:0] s_282;
  wire [0:0] s_283;
  wire [0:0] s_284;
  wire [0:0] s_285;
  wire [0:0] s_286;
  wire [0:0] s_287;
  wire [2:0] s_288;
  wire [0:0] s_289;
  wire [0:0] s_290;
  wire [1:0] s_291;
  wire [1:0] s_292;
  wire [1:0] s_293;
  wire [3:0] s_294;
  wire [0:0] s_295;
  wire [0:0] s_296;
  wire [2:0] s_297;
  wire [2:0] s_298;
  wire [2:0] s_299;
  wire [0:0] s_300;
  wire [4:0] s_301;
  wire [0:0] s_302;
  wire [0:0] s_303;
  wire [3:0] s_304;
  wire [0:0] s_305;
  wire [0:0] s_306;
  wire [2:0] s_307;
  wire [0:0] s_308;
  wire [0:0] s_309;
  wire [1:0] s_310;
  wire [0:0] s_311;
  wire [0:0] s_312;
  wire [0:0] s_313;
  wire [1:0] s_314;
  wire [3:0] s_315;
  wire [7:0] s_316;
  wire [15:0] s_317;
  wire [0:0] s_318;
  wire [0:0] s_319;
  wire [0:0] s_320;
  wire [0:0] s_321;
  wire [0:0] s_322;
  wire [0:0] s_323;
  wire [0:0] s_324;
  wire [1:0] s_325;
  wire [0:0] s_326;
  wire [0:0] s_327;
  wire [0:0] s_328;
  wire [1:0] s_329;
  wire [0:0] s_330;
  wire [0:0] s_331;
  wire [0:0] s_332;
  wire [0:0] s_333;
  wire [0:0] s_334;
  wire [0:0] s_335;
  wire [1:0] s_336;
  wire [0:0] s_337;
  wire [0:0] s_338;
  wire [0:0] s_339;
  wire [0:0] s_340;
  wire [0:0] s_341;
  wire [0:0] s_342;
  wire [2:0] s_343;
  wire [0:0] s_344;
  wire [0:0] s_345;
  wire [1:0] s_346;
  wire [0:0] s_347;
  wire [0:0] s_348;
  wire [0:0] s_349;
  wire [1:0] s_350;
  wire [3:0] s_351;
  wire [0:0] s_352;
  wire [0:0] s_353;
  wire [0:0] s_354;
  wire [0:0] s_355;
  wire [0:0] s_356;
  wire [0:0] s_357;
  wire [0:0] s_358;
  wire [1:0] s_359;
  wire [0:0] s_360;
  wire [0:0] s_361;
  wire [0:0] s_362;
  wire [1:0] s_363;
  wire [0:0] s_364;
  wire [0:0] s_365;
  wire [0:0] s_366;
  wire [0:0] s_367;
  wire [0:0] s_368;
  wire [0:0] s_369;
  wire [1:0] s_370;
  wire [0:0] s_371;
  wire [0:0] s_372;
  wire [0:0] s_373;
  wire [0:0] s_374;
  wire [0:0] s_375;
  wire [2:0] s_376;
  wire [0:0] s_377;
  wire [0:0] s_378;
  wire [1:0] s_379;
  wire [1:0] s_380;
  wire [1:0] s_381;
  wire [0:0] s_382;
  wire [3:0] s_383;
  wire [0:0] s_384;
  wire [0:0] s_385;
  wire [2:0] s_386;
  wire [0:0] s_387;
  wire [0:0] s_388;
  wire [1:0] s_389;
  wire [0:0] s_390;
  wire [0:0] s_391;
  wire [0:0] s_392;
  wire [1:0] s_393;
  wire [3:0] s_394;
  wire [7:0] s_395;
  wire [0:0] s_396;
  wire [0:0] s_397;
  wire [0:0] s_398;
  wire [0:0] s_399;
  wire [0:0] s_400;
  wire [0:0] s_401;
  wire [0:0] s_402;
  wire [1:0] s_403;
  wire [0:0] s_404;
  wire [0:0] s_405;
  wire [0:0] s_406;
  wire [1:0] s_407;
  wire [0:0] s_408;
  wire [0:0] s_409;
  wire [0:0] s_410;
  wire [0:0] s_411;
  wire [0:0] s_412;
  wire [0:0] s_413;
  wire [1:0] s_414;
  wire [0:0] s_415;
  wire [0:0] s_416;
  wire [0:0] s_417;
  wire [0:0] s_418;
  wire [0:0] s_419;
  wire [0:0] s_420;
  wire [2:0] s_421;
  wire [0:0] s_422;
  wire [0:0] s_423;
  wire [1:0] s_424;
  wire [0:0] s_425;
  wire [0:0] s_426;
  wire [0:0] s_427;
  wire [1:0] s_428;
  wire [3:0] s_429;
  wire [0:0] s_430;
  wire [0:0] s_431;
  wire [0:0] s_432;
  wire [0:0] s_433;
  wire [0:0] s_434;
  wire [0:0] s_435;
  wire [0:0] s_436;
  wire [1:0] s_437;
  wire [0:0] s_438;
  wire [0:0] s_439;
  wire [0:0] s_440;
  wire [1:0] s_441;
  wire [0:0] s_442;
  wire [0:0] s_443;
  wire [0:0] s_444;
  wire [0:0] s_445;
  wire [0:0] s_446;
  wire [0:0] s_447;
  wire [1:0] s_448;
  wire [0:0] s_449;
  wire [0:0] s_450;
  wire [0:0] s_451;
  wire [0:0] s_452;
  wire [0:0] s_453;
  wire [2:0] s_454;
  wire [0:0] s_455;
  wire [0:0] s_456;
  wire [1:0] s_457;
  wire [1:0] s_458;
  wire [1:0] s_459;
  wire [3:0] s_460;
  wire [0:0] s_461;
  wire [0:0] s_462;
  wire [2:0] s_463;
  wire [2:0] s_464;
  wire [2:0] s_465;
  wire [4:0] s_466;
  wire [0:0] s_467;
  wire [0:0] s_468;
  wire [3:0] s_469;
  wire [3:0] s_470;
  wire [3:0] s_471;
  wire [0:0] s_472;
  wire [5:0] s_473;
  wire [0:0] s_474;
  wire [0:0] s_475;
  wire [4:0] s_476;
  wire [0:0] s_477;
  wire [0:0] s_478;
  wire [3:0] s_479;
  wire [0:0] s_480;
  wire [0:0] s_481;
  wire [2:0] s_482;
  wire [0:0] s_483;
  wire [0:0] s_484;
  wire [1:0] s_485;
  wire [0:0] s_486;
  wire [0:0] s_487;
  wire [0:0] s_488;
  wire [1:0] s_489;
  wire [3:0] s_490;
  wire [7:0] s_491;
  wire [15:0] s_492;
  wire [31:0] s_493;
  wire [0:0] s_494;
  wire [0:0] s_495;
  wire [0:0] s_496;
  wire [0:0] s_497;
  wire [0:0] s_498;
  wire [0:0] s_499;
  wire [0:0] s_500;
  wire [1:0] s_501;
  wire [0:0] s_502;
  wire [0:0] s_503;
  wire [0:0] s_504;
  wire [1:0] s_505;
  wire [0:0] s_506;
  wire [0:0] s_507;
  wire [0:0] s_508;
  wire [0:0] s_509;
  wire [0:0] s_510;
  wire [0:0] s_511;
  wire [1:0] s_512;
  wire [0:0] s_513;
  wire [0:0] s_514;
  wire [0:0] s_515;
  wire [0:0] s_516;
  wire [0:0] s_517;
  wire [0:0] s_518;
  wire [2:0] s_519;
  wire [0:0] s_520;
  wire [0:0] s_521;
  wire [1:0] s_522;
  wire [0:0] s_523;
  wire [0:0] s_524;
  wire [0:0] s_525;
  wire [1:0] s_526;
  wire [3:0] s_527;
  wire [0:0] s_528;
  wire [0:0] s_529;
  wire [0:0] s_530;
  wire [0:0] s_531;
  wire [0:0] s_532;
  wire [0:0] s_533;
  wire [0:0] s_534;
  wire [1:0] s_535;
  wire [0:0] s_536;
  wire [0:0] s_537;
  wire [0:0] s_538;
  wire [1:0] s_539;
  wire [0:0] s_540;
  wire [0:0] s_541;
  wire [0:0] s_542;
  wire [0:0] s_543;
  wire [0:0] s_544;
  wire [0:0] s_545;
  wire [1:0] s_546;
  wire [0:0] s_547;
  wire [0:0] s_548;
  wire [0:0] s_549;
  wire [0:0] s_550;
  wire [0:0] s_551;
  wire [2:0] s_552;
  wire [0:0] s_553;
  wire [0:0] s_554;
  wire [1:0] s_555;
  wire [1:0] s_556;
  wire [1:0] s_557;
  wire [0:0] s_558;
  wire [3:0] s_559;
  wire [0:0] s_560;
  wire [0:0] s_561;
  wire [2:0] s_562;
  wire [0:0] s_563;
  wire [0:0] s_564;
  wire [1:0] s_565;
  wire [0:0] s_566;
  wire [0:0] s_567;
  wire [0:0] s_568;
  wire [1:0] s_569;
  wire [3:0] s_570;
  wire [7:0] s_571;
  wire [0:0] s_572;
  wire [0:0] s_573;
  wire [0:0] s_574;
  wire [0:0] s_575;
  wire [0:0] s_576;
  wire [0:0] s_577;
  wire [0:0] s_578;
  wire [1:0] s_579;
  wire [0:0] s_580;
  wire [0:0] s_581;
  wire [0:0] s_582;
  wire [1:0] s_583;
  wire [0:0] s_584;
  wire [0:0] s_585;
  wire [0:0] s_586;
  wire [0:0] s_587;
  wire [0:0] s_588;
  wire [0:0] s_589;
  wire [1:0] s_590;
  wire [0:0] s_591;
  wire [0:0] s_592;
  wire [0:0] s_593;
  wire [0:0] s_594;
  wire [0:0] s_595;
  wire [0:0] s_596;
  wire [2:0] s_597;
  wire [0:0] s_598;
  wire [0:0] s_599;
  wire [1:0] s_600;
  wire [0:0] s_601;
  wire [0:0] s_602;
  wire [0:0] s_603;
  wire [1:0] s_604;
  wire [3:0] s_605;
  wire [0:0] s_606;
  wire [0:0] s_607;
  wire [0:0] s_608;
  wire [0:0] s_609;
  wire [0:0] s_610;
  wire [0:0] s_611;
  wire [0:0] s_612;
  wire [1:0] s_613;
  wire [0:0] s_614;
  wire [0:0] s_615;
  wire [0:0] s_616;
  wire [1:0] s_617;
  wire [0:0] s_618;
  wire [0:0] s_619;
  wire [0:0] s_620;
  wire [0:0] s_621;
  wire [0:0] s_622;
  wire [0:0] s_623;
  wire [1:0] s_624;
  wire [0:0] s_625;
  wire [0:0] s_626;
  wire [0:0] s_627;
  wire [0:0] s_628;
  wire [0:0] s_629;
  wire [2:0] s_630;
  wire [0:0] s_631;
  wire [0:0] s_632;
  wire [1:0] s_633;
  wire [1:0] s_634;
  wire [1:0] s_635;
  wire [3:0] s_636;
  wire [0:0] s_637;
  wire [0:0] s_638;
  wire [2:0] s_639;
  wire [2:0] s_640;
  wire [2:0] s_641;
  wire [0:0] s_642;
  wire [4:0] s_643;
  wire [0:0] s_644;
  wire [0:0] s_645;
  wire [3:0] s_646;
  wire [0:0] s_647;
  wire [0:0] s_648;
  wire [2:0] s_649;
  wire [0:0] s_650;
  wire [0:0] s_651;
  wire [1:0] s_652;
  wire [0:0] s_653;
  wire [0:0] s_654;
  wire [0:0] s_655;
  wire [1:0] s_656;
  wire [3:0] s_657;
  wire [7:0] s_658;
  wire [15:0] s_659;
  wire [0:0] s_660;
  wire [0:0] s_661;
  wire [0:0] s_662;
  wire [0:0] s_663;
  wire [0:0] s_664;
  wire [0:0] s_665;
  wire [0:0] s_666;
  wire [1:0] s_667;
  wire [0:0] s_668;
  wire [0:0] s_669;
  wire [0:0] s_670;
  wire [1:0] s_671;
  wire [0:0] s_672;
  wire [0:0] s_673;
  wire [0:0] s_674;
  wire [0:0] s_675;
  wire [0:0] s_676;
  wire [0:0] s_677;
  wire [1:0] s_678;
  wire [0:0] s_679;
  wire [0:0] s_680;
  wire [0:0] s_681;
  wire [0:0] s_682;
  wire [0:0] s_683;
  wire [0:0] s_684;
  wire [2:0] s_685;
  wire [0:0] s_686;
  wire [0:0] s_687;
  wire [1:0] s_688;
  wire [0:0] s_689;
  wire [0:0] s_690;
  wire [0:0] s_691;
  wire [1:0] s_692;
  wire [3:0] s_693;
  wire [0:0] s_694;
  wire [0:0] s_695;
  wire [0:0] s_696;
  wire [0:0] s_697;
  wire [0:0] s_698;
  wire [0:0] s_699;
  wire [0:0] s_700;
  wire [1:0] s_701;
  wire [0:0] s_702;
  wire [0:0] s_703;
  wire [0:0] s_704;
  wire [1:0] s_705;
  wire [0:0] s_706;
  wire [0:0] s_707;
  wire [0:0] s_708;
  wire [0:0] s_709;
  wire [0:0] s_710;
  wire [0:0] s_711;
  wire [1:0] s_712;
  wire [0:0] s_713;
  wire [0:0] s_714;
  wire [0:0] s_715;
  wire [0:0] s_716;
  wire [0:0] s_717;
  wire [2:0] s_718;
  wire [0:0] s_719;
  wire [0:0] s_720;
  wire [1:0] s_721;
  wire [1:0] s_722;
  wire [1:0] s_723;
  wire [0:0] s_724;
  wire [3:0] s_725;
  wire [0:0] s_726;
  wire [0:0] s_727;
  wire [2:0] s_728;
  wire [0:0] s_729;
  wire [0:0] s_730;
  wire [1:0] s_731;
  wire [0:0] s_732;
  wire [0:0] s_733;
  wire [0:0] s_734;
  wire [1:0] s_735;
  wire [3:0] s_736;
  wire [7:0] s_737;
  wire [0:0] s_738;
  wire [0:0] s_739;
  wire [0:0] s_740;
  wire [0:0] s_741;
  wire [0:0] s_742;
  wire [0:0] s_743;
  wire [0:0] s_744;
  wire [1:0] s_745;
  wire [0:0] s_746;
  wire [0:0] s_747;
  wire [0:0] s_748;
  wire [1:0] s_749;
  wire [0:0] s_750;
  wire [0:0] s_751;
  wire [0:0] s_752;
  wire [0:0] s_753;
  wire [0:0] s_754;
  wire [0:0] s_755;
  wire [1:0] s_756;
  wire [0:0] s_757;
  wire [0:0] s_758;
  wire [0:0] s_759;
  wire [0:0] s_760;
  wire [0:0] s_761;
  wire [0:0] s_762;
  wire [2:0] s_763;
  wire [0:0] s_764;
  wire [0:0] s_765;
  wire [1:0] s_766;
  wire [0:0] s_767;
  wire [0:0] s_768;
  wire [0:0] s_769;
  wire [1:0] s_770;
  wire [3:0] s_771;
  wire [0:0] s_772;
  wire [0:0] s_773;
  wire [0:0] s_774;
  wire [0:0] s_775;
  wire [0:0] s_776;
  wire [0:0] s_777;
  wire [0:0] s_778;
  wire [1:0] s_779;
  wire [0:0] s_780;
  wire [0:0] s_781;
  wire [0:0] s_782;
  wire [1:0] s_783;
  wire [0:0] s_784;
  wire [0:0] s_785;
  wire [0:0] s_786;
  wire [0:0] s_787;
  wire [0:0] s_788;
  wire [0:0] s_789;
  wire [1:0] s_790;
  wire [0:0] s_791;
  wire [0:0] s_792;
  wire [0:0] s_793;
  wire [0:0] s_794;
  wire [0:0] s_795;
  wire [2:0] s_796;
  wire [0:0] s_797;
  wire [0:0] s_798;
  wire [1:0] s_799;
  wire [1:0] s_800;
  wire [1:0] s_801;
  wire [3:0] s_802;
  wire [0:0] s_803;
  wire [0:0] s_804;
  wire [2:0] s_805;
  wire [2:0] s_806;
  wire [2:0] s_807;
  wire [4:0] s_808;
  wire [0:0] s_809;
  wire [0:0] s_810;
  wire [3:0] s_811;
  wire [3:0] s_812;
  wire [3:0] s_813;
  wire [5:0] s_814;
  wire [0:0] s_815;
  wire [0:0] s_816;
  wire [4:0] s_817;
  wire [4:0] s_818;
  wire [4:0] s_819;
  wire [11:0] s_820;
  wire [11:0] s_821;
  wire [11:0] s_822;
  wire [11:0] s_823;
  wire [11:0] s_824;
  wire [11:0] s_825;
  wire [0:0] s_826;
  wire [11:0] s_827;
  wire [0:0] s_828;
  wire [11:0] s_829;
  wire [11:0] s_830;
  wire [0:0] s_831;
  wire [52:0] s_832;
  wire [0:0] s_833;
  wire [0:0] s_834;
  wire [0:0] s_835;
  wire [0:0] s_836;
  wire [0:0] s_837;
  wire [0:0] s_838;
  wire [0:0] s_839;
  wire [0:0] s_840;
  wire [0:0] s_841;
  wire [0:0] s_842;
  wire [0:0] s_843;
  wire [0:0] s_844;
  wire [0:0] s_845;
  wire [52:0] s_846;
  wire [0:0] s_847;
  wire [63:0] s_848;
  wire [11:0] s_849;
  wire [0:0] s_850;
  wire [10:0] s_851;
  wire [10:0] s_852;
  wire [11:0] s_853;
  wire [11:0] s_854;
  wire [11:0] s_855;
  wire [11:0] s_856;
  wire [11:0] s_857;
  wire [11:0] s_858;
  wire [9:0] s_859;
  wire [51:0] s_860;
  wire [0:0] s_861;
  wire [0:0] s_862;
  wire [10:0] s_863;
  wire [0:0] s_864;
  wire [0:0] s_865;
  wire [0:0] s_866;
  wire [52:0] s_867;
  wire [0:0] s_868;
  wire [0:0] s_869;
  wire [0:0] s_870;
  wire [10:0] s_871;
  wire [0:0] s_872;
  wire [0:0] s_873;
  wire [0:0] s_874;
  wire [0:0] s_875;
  wire [0:0] s_876;
  wire [0:0] s_877;
  wire [0:0] s_878;
  wire [10:0] s_879;
  wire [0:0] s_880;
  wire [51:0] s_881;
  wire [0:0] s_882;
  wire [0:0] s_883;
  wire [10:0] s_884;
  wire [0:0] s_885;
  wire [51:0] s_886;
  wire [0:0] s_887;

  assign s_0 = s_874?s_1:s_85;
  dq #(64, 5) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_84};
  assign s_3 = s_72?s_4:s_5;
  assign s_4 = 1'd0;
  dq #(1, 2) dq_s_5 (clk, s_5, s_6);
  assign s_6 = s_45?s_7:s_44;
  assign s_7 = s_12?s_8:s_10;
  assign s_8 = s_9[63];
  assign s_9 = double_add_a;
  assign s_10 = s_11[63];
  assign s_11 = double_add_b;
  assign s_12 = s_13 & s_37;
  assign s_13 = s_14 | s_31;
  assign s_14 = $signed(s_15) > $signed(s_23);
  assign s_15 = $signed(s_16);
  assign s_16 = s_21?s_17:s_18;
  assign s_17 = -11'd1022;
  assign s_18 = s_19 - s_20;
  assign s_19 = s_9[62:52];
  assign s_20 = 10'd1023;
  assign s_21 = s_18 == s_22;
  assign s_22 = -11'd1023;
  assign s_23 = $signed(s_24);
  assign s_24 = s_29?s_25:s_26;
  assign s_25 = -11'd1022;
  assign s_26 = s_27 - s_28;
  assign s_27 = s_11[62:52];
  assign s_28 = 10'd1023;
  assign s_29 = s_26 == s_30;
  assign s_30 = -11'd1023;
  assign s_31 = s_32 & s_34;
  assign s_32 = s_18 == s_33;
  assign s_33 = 11'd1024;
  assign s_34 = s_35 == s_36;
  assign s_35 = s_9[51:0];
  assign s_36 = 52'd0;
  assign s_37 = ~s_38;
  assign s_38 = s_39 & s_41;
  assign s_39 = s_26 == s_40;
  assign s_40 = 11'd1024;
  assign s_41 = s_42 == s_43;
  assign s_42 = s_11[51:0];
  assign s_43 = 52'd0;
  assign s_44 = s_12?s_10:s_8;
  assign s_45 = s_46 >= s_58;
  assign s_46 = s_47 << s_57;
  assign s_47 = s_48;
  assign s_48 = s_12?s_49:s_53;
  assign s_49 = {s_50,s_35};
  assign s_50 = s_21?s_51:s_52;
  assign s_51 = 1'd0;
  assign s_52 = 1'd1;
  assign s_53 = {s_54,s_42};
  assign s_54 = s_29?s_55:s_56;
  assign s_55 = 1'd0;
  assign s_56 = 1'd1;
  assign s_57 = 2'd3;
  assign s_58 = s_59 | s_67;
  assign s_59 = s_60 >> s_64;
  assign s_60 = s_61 << s_63;
  assign s_61 = s_62;
  assign s_62 = s_12?s_53:s_49;
  assign s_63 = 2'd3;
  assign s_64 = s_65 - s_66;
  assign s_65 = s_12?s_15:s_23;
  assign s_66 = s_12?s_23:s_15;
  assign s_67 = s_68 != s_71;
  assign s_68 = s_60 << s_69;
  assign s_69 = s_70 - s_64;
  assign s_70 = 57'd57;
  assign s_71 = 1'd0;
  assign s_72 = s_73 == s_83;
  dq #(57, 1) dq_s_73 (clk, s_73, s_74);
  assign s_74 = s_75 + s_77;
  dq #(57, 1) dq_s_75 (clk, s_75, s_76);
  assign s_76 = s_45?s_46:s_58;
  dq #(57, 1) dq_s_77 (clk, s_77, s_78);
  assign s_78 = s_82?s_79:s_80;
  assign s_79 = s_45?s_58:s_46;
  assign s_80 = s_81 - s_79;
  assign s_81 = 57'd0;
  assign s_82 = s_8 == s_10;
  assign s_83 = 1'd0;
  assign s_84 = 63'd9221120237041090560;
  assign s_85 = s_868?s_86:s_89;
  dq #(64, 5) dq_s_86 (clk, s_86, s_87);
  assign s_87 = {s_3,s_88};
  assign s_88 = 63'd9218868437227405312;
  assign s_89 = s_866?s_90:s_93;
  dq #(64, 5) dq_s_90 (clk, s_90, s_91);
  assign s_91 = {s_3,s_92};
  assign s_92 = 63'd0;
  assign s_93 = s_861?s_94:s_848;
  assign s_94 = {s_95,s_98};
  dq #(12, 5) dq_s_95 (clk, s_95, s_96);
  assign s_96 = {s_3,s_97};
  assign s_97 = 11'd0;
  assign s_98 = s_99[51:0];
  dq #(53, 1) dq_s_99 (clk, s_99, s_100);
  assign s_100 = s_847?s_101:s_846;
  assign s_101 = s_102[53:1];
  assign s_102 = s_833?s_103:s_832;
  dq #(54, 1) dq_s_103 (clk, s_103, s_104);
  assign s_104 = s_105 + s_831;
  assign s_105 = s_106;
  assign s_106 = s_107[56:4];
  dq #(57, 1) dq_s_107 (clk, s_107, s_108);
  assign s_108 = s_109 << s_111;
  dq #(57, 2) dq_s_109 (clk, s_109, s_110);
  dq #(57, 1) dq_s_110 (clk, s_110, s_74);
  dq #(12, 1) dq_s_111 (clk, s_111, s_112);
  assign s_112 = s_828?s_113:s_820;
  dq #(7, 1) dq_s_113 (clk, s_113, s_114);
  assign s_114 = {s_115,s_814};
  assign s_115 = s_116 & s_472;
  assign s_116 = s_117[5];
  assign s_117 = {s_118,s_466};
  assign s_118 = s_119 & s_300;
  assign s_119 = s_120[4];
  assign s_120 = {s_121,s_294};
  assign s_121 = s_122 & s_216;
  assign s_122 = s_123[3];
  assign s_123 = {s_124,s_210};
  assign s_124 = s_125 & s_176;
  assign s_125 = s_126[2];
  assign s_126 = {s_127,s_170};
  assign s_127 = s_128 & s_158;
  assign s_128 = s_129[1];
  assign s_129 = {s_130,s_154};
  assign s_130 = s_131 & s_152;
  assign s_131 = ~s_132;
  assign s_132 = s_133[1];
  assign s_133 = s_134[3:2];
  assign s_134 = s_135[7:4];
  assign s_135 = s_136[15:8];
  assign s_136 = s_137[31:16];
  assign s_137 = s_138[63:32];
  assign s_138 = {s_139,s_151};
  assign s_139 = {s_140,s_150};
  assign s_140 = {s_141,s_149};
  assign s_141 = {s_142,s_148};
  assign s_142 = {s_143,s_147};
  assign s_143 = {s_144,s_146};
  assign s_144 = {s_110,s_145};
  assign s_145 = 1'd1;
  assign s_146 = 1'd1;
  assign s_147 = 1'd1;
  assign s_148 = 1'd1;
  assign s_149 = 1'd1;
  assign s_150 = 1'd1;
  assign s_151 = 1'd1;
  assign s_152 = ~s_153;
  assign s_153 = s_133[0];
  assign s_154 = s_155 & s_157;
  assign s_155 = ~s_156;
  assign s_156 = s_133[1];
  assign s_157 = s_133[0];
  assign s_158 = s_159[1];
  assign s_159 = {s_160,s_166};
  assign s_160 = s_161 & s_164;
  assign s_161 = ~s_162;
  assign s_162 = s_163[1];
  assign s_163 = s_134[1:0];
  assign s_164 = ~s_165;
  assign s_165 = s_163[0];
  assign s_166 = s_167 & s_169;
  assign s_167 = ~s_168;
  assign s_168 = s_163[1];
  assign s_169 = s_163[0];
  assign s_170 = {s_171,s_173};
  assign s_171 = s_128 & s_172;
  assign s_172 = ~s_158;
  assign s_173 = s_128?s_174:s_175;
  assign s_174 = s_159[0:0];
  assign s_175 = s_129[0:0];
  assign s_176 = s_177[2];
  assign s_177 = {s_178,s_204};
  assign s_178 = s_179 & s_192;
  assign s_179 = s_180[1];
  assign s_180 = {s_181,s_188};
  assign s_181 = s_182 & s_186;
  assign s_182 = ~s_183;
  assign s_183 = s_184[1];
  assign s_184 = s_185[3:2];
  assign s_185 = s_135[3:0];
  assign s_186 = ~s_187;
  assign s_187 = s_184[0];
  assign s_188 = s_189 & s_191;
  assign s_189 = ~s_190;
  assign s_190 = s_184[1];
  assign s_191 = s_184[0];
  assign s_192 = s_193[1];
  assign s_193 = {s_194,s_200};
  assign s_194 = s_195 & s_198;
  assign s_195 = ~s_196;
  assign s_196 = s_197[1];
  assign s_197 = s_185[1:0];
  assign s_198 = ~s_199;
  assign s_199 = s_197[0];
  assign s_200 = s_201 & s_203;
  assign s_201 = ~s_202;
  assign s_202 = s_197[1];
  assign s_203 = s_197[0];
  assign s_204 = {s_205,s_207};
  assign s_205 = s_179 & s_206;
  assign s_206 = ~s_192;
  assign s_207 = s_179?s_208:s_209;
  assign s_208 = s_193[0:0];
  assign s_209 = s_180[0:0];
  assign s_210 = {s_211,s_213};
  assign s_211 = s_125 & s_212;
  assign s_212 = ~s_176;
  assign s_213 = s_125?s_214:s_215;
  assign s_214 = s_177[1:0];
  assign s_215 = s_126[1:0];
  assign s_216 = s_217[3];
  assign s_217 = {s_218,s_288};
  assign s_218 = s_219 & s_254;
  assign s_219 = s_220[2];
  assign s_220 = {s_221,s_248};
  assign s_221 = s_222 & s_236;
  assign s_222 = s_223[1];
  assign s_223 = {s_224,s_232};
  assign s_224 = s_225 & s_230;
  assign s_225 = ~s_226;
  assign s_226 = s_227[1];
  assign s_227 = s_228[3:2];
  assign s_228 = s_229[7:4];
  assign s_229 = s_136[7:0];
  assign s_230 = ~s_231;
  assign s_231 = s_227[0];
  assign s_232 = s_233 & s_235;
  assign s_233 = ~s_234;
  assign s_234 = s_227[1];
  assign s_235 = s_227[0];
  assign s_236 = s_237[1];
  assign s_237 = {s_238,s_244};
  assign s_238 = s_239 & s_242;
  assign s_239 = ~s_240;
  assign s_240 = s_241[1];
  assign s_241 = s_228[1:0];
  assign s_242 = ~s_243;
  assign s_243 = s_241[0];
  assign s_244 = s_245 & s_247;
  assign s_245 = ~s_246;
  assign s_246 = s_241[1];
  assign s_247 = s_241[0];
  assign s_248 = {s_249,s_251};
  assign s_249 = s_222 & s_250;
  assign s_250 = ~s_236;
  assign s_251 = s_222?s_252:s_253;
  assign s_252 = s_237[0:0];
  assign s_253 = s_223[0:0];
  assign s_254 = s_255[2];
  assign s_255 = {s_256,s_282};
  assign s_256 = s_257 & s_270;
  assign s_257 = s_258[1];
  assign s_258 = {s_259,s_266};
  assign s_259 = s_260 & s_264;
  assign s_260 = ~s_261;
  assign s_261 = s_262[1];
  assign s_262 = s_263[3:2];
  assign s_263 = s_229[3:0];
  assign s_264 = ~s_265;
  assign s_265 = s_262[0];
  assign s_266 = s_267 & s_269;
  assign s_267 = ~s_268;
  assign s_268 = s_262[1];
  assign s_269 = s_262[0];
  assign s_270 = s_271[1];
  assign s_271 = {s_272,s_278};
  assign s_272 = s_273 & s_276;
  assign s_273 = ~s_274;
  assign s_274 = s_275[1];
  assign s_275 = s_263[1:0];
  assign s_276 = ~s_277;
  assign s_277 = s_275[0];
  assign s_278 = s_279 & s_281;
  assign s_279 = ~s_280;
  assign s_280 = s_275[1];
  assign s_281 = s_275[0];
  assign s_282 = {s_283,s_285};
  assign s_283 = s_257 & s_284;
  assign s_284 = ~s_270;
  assign s_285 = s_257?s_286:s_287;
  assign s_286 = s_271[0:0];
  assign s_287 = s_258[0:0];
  assign s_288 = {s_289,s_291};
  assign s_289 = s_219 & s_290;
  assign s_290 = ~s_254;
  assign s_291 = s_219?s_292:s_293;
  assign s_292 = s_255[1:0];
  assign s_293 = s_220[1:0];
  assign s_294 = {s_295,s_297};
  assign s_295 = s_122 & s_296;
  assign s_296 = ~s_216;
  assign s_297 = s_122?s_298:s_299;
  assign s_298 = s_217[2:0];
  assign s_299 = s_123[2:0];
  assign s_300 = s_301[4];
  assign s_301 = {s_302,s_460};
  assign s_302 = s_303 & s_382;
  assign s_303 = s_304[3];
  assign s_304 = {s_305,s_376};
  assign s_305 = s_306 & s_342;
  assign s_306 = s_307[2];
  assign s_307 = {s_308,s_336};
  assign s_308 = s_309 & s_324;
  assign s_309 = s_310[1];
  assign s_310 = {s_311,s_320};
  assign s_311 = s_312 & s_318;
  assign s_312 = ~s_313;
  assign s_313 = s_314[1];
  assign s_314 = s_315[3:2];
  assign s_315 = s_316[7:4];
  assign s_316 = s_317[15:8];
  assign s_317 = s_137[15:0];
  assign s_318 = ~s_319;
  assign s_319 = s_314[0];
  assign s_320 = s_321 & s_323;
  assign s_321 = ~s_322;
  assign s_322 = s_314[1];
  assign s_323 = s_314[0];
  assign s_324 = s_325[1];
  assign s_325 = {s_326,s_332};
  assign s_326 = s_327 & s_330;
  assign s_327 = ~s_328;
  assign s_328 = s_329[1];
  assign s_329 = s_315[1:0];
  assign s_330 = ~s_331;
  assign s_331 = s_329[0];
  assign s_332 = s_333 & s_335;
  assign s_333 = ~s_334;
  assign s_334 = s_329[1];
  assign s_335 = s_329[0];
  assign s_336 = {s_337,s_339};
  assign s_337 = s_309 & s_338;
  assign s_338 = ~s_324;
  assign s_339 = s_309?s_340:s_341;
  assign s_340 = s_325[0:0];
  assign s_341 = s_310[0:0];
  assign s_342 = s_343[2];
  assign s_343 = {s_344,s_370};
  assign s_344 = s_345 & s_358;
  assign s_345 = s_346[1];
  assign s_346 = {s_347,s_354};
  assign s_347 = s_348 & s_352;
  assign s_348 = ~s_349;
  assign s_349 = s_350[1];
  assign s_350 = s_351[3:2];
  assign s_351 = s_316[3:0];
  assign s_352 = ~s_353;
  assign s_353 = s_350[0];
  assign s_354 = s_355 & s_357;
  assign s_355 = ~s_356;
  assign s_356 = s_350[1];
  assign s_357 = s_350[0];
  assign s_358 = s_359[1];
  assign s_359 = {s_360,s_366};
  assign s_360 = s_361 & s_364;
  assign s_361 = ~s_362;
  assign s_362 = s_363[1];
  assign s_363 = s_351[1:0];
  assign s_364 = ~s_365;
  assign s_365 = s_363[0];
  assign s_366 = s_367 & s_369;
  assign s_367 = ~s_368;
  assign s_368 = s_363[1];
  assign s_369 = s_363[0];
  assign s_370 = {s_371,s_373};
  assign s_371 = s_345 & s_372;
  assign s_372 = ~s_358;
  assign s_373 = s_345?s_374:s_375;
  assign s_374 = s_359[0:0];
  assign s_375 = s_346[0:0];
  assign s_376 = {s_377,s_379};
  assign s_377 = s_306 & s_378;
  assign s_378 = ~s_342;
  assign s_379 = s_306?s_380:s_381;
  assign s_380 = s_343[1:0];
  assign s_381 = s_307[1:0];
  assign s_382 = s_383[3];
  assign s_383 = {s_384,s_454};
  assign s_384 = s_385 & s_420;
  assign s_385 = s_386[2];
  assign s_386 = {s_387,s_414};
  assign s_387 = s_388 & s_402;
  assign s_388 = s_389[1];
  assign s_389 = {s_390,s_398};
  assign s_390 = s_391 & s_396;
  assign s_391 = ~s_392;
  assign s_392 = s_393[1];
  assign s_393 = s_394[3:2];
  assign s_394 = s_395[7:4];
  assign s_395 = s_317[7:0];
  assign s_396 = ~s_397;
  assign s_397 = s_393[0];
  assign s_398 = s_399 & s_401;
  assign s_399 = ~s_400;
  assign s_400 = s_393[1];
  assign s_401 = s_393[0];
  assign s_402 = s_403[1];
  assign s_403 = {s_404,s_410};
  assign s_404 = s_405 & s_408;
  assign s_405 = ~s_406;
  assign s_406 = s_407[1];
  assign s_407 = s_394[1:0];
  assign s_408 = ~s_409;
  assign s_409 = s_407[0];
  assign s_410 = s_411 & s_413;
  assign s_411 = ~s_412;
  assign s_412 = s_407[1];
  assign s_413 = s_407[0];
  assign s_414 = {s_415,s_417};
  assign s_415 = s_388 & s_416;
  assign s_416 = ~s_402;
  assign s_417 = s_388?s_418:s_419;
  assign s_418 = s_403[0:0];
  assign s_419 = s_389[0:0];
  assign s_420 = s_421[2];
  assign s_421 = {s_422,s_448};
  assign s_422 = s_423 & s_436;
  assign s_423 = s_424[1];
  assign s_424 = {s_425,s_432};
  assign s_425 = s_426 & s_430;
  assign s_426 = ~s_427;
  assign s_427 = s_428[1];
  assign s_428 = s_429[3:2];
  assign s_429 = s_395[3:0];
  assign s_430 = ~s_431;
  assign s_431 = s_428[0];
  assign s_432 = s_433 & s_435;
  assign s_433 = ~s_434;
  assign s_434 = s_428[1];
  assign s_435 = s_428[0];
  assign s_436 = s_437[1];
  assign s_437 = {s_438,s_444};
  assign s_438 = s_439 & s_442;
  assign s_439 = ~s_440;
  assign s_440 = s_441[1];
  assign s_441 = s_429[1:0];
  assign s_442 = ~s_443;
  assign s_443 = s_441[0];
  assign s_444 = s_445 & s_447;
  assign s_445 = ~s_446;
  assign s_446 = s_441[1];
  assign s_447 = s_441[0];
  assign s_448 = {s_449,s_451};
  assign s_449 = s_423 & s_450;
  assign s_450 = ~s_436;
  assign s_451 = s_423?s_452:s_453;
  assign s_452 = s_437[0:0];
  assign s_453 = s_424[0:0];
  assign s_454 = {s_455,s_457};
  assign s_455 = s_385 & s_456;
  assign s_456 = ~s_420;
  assign s_457 = s_385?s_458:s_459;
  assign s_458 = s_421[1:0];
  assign s_459 = s_386[1:0];
  assign s_460 = {s_461,s_463};
  assign s_461 = s_303 & s_462;
  assign s_462 = ~s_382;
  assign s_463 = s_303?s_464:s_465;
  assign s_464 = s_383[2:0];
  assign s_465 = s_304[2:0];
  assign s_466 = {s_467,s_469};
  assign s_467 = s_119 & s_468;
  assign s_468 = ~s_300;
  assign s_469 = s_119?s_470:s_471;
  assign s_470 = s_301[3:0];
  assign s_471 = s_120[3:0];
  assign s_472 = s_473[5];
  assign s_473 = {s_474,s_808};
  assign s_474 = s_475 & s_642;
  assign s_475 = s_476[4];
  assign s_476 = {s_477,s_636};
  assign s_477 = s_478 & s_558;
  assign s_478 = s_479[3];
  assign s_479 = {s_480,s_552};
  assign s_480 = s_481 & s_518;
  assign s_481 = s_482[2];
  assign s_482 = {s_483,s_512};
  assign s_483 = s_484 & s_500;
  assign s_484 = s_485[1];
  assign s_485 = {s_486,s_496};
  assign s_486 = s_487 & s_494;
  assign s_487 = ~s_488;
  assign s_488 = s_489[1];
  assign s_489 = s_490[3:2];
  assign s_490 = s_491[7:4];
  assign s_491 = s_492[15:8];
  assign s_492 = s_493[31:16];
  assign s_493 = s_138[31:0];
  assign s_494 = ~s_495;
  assign s_495 = s_489[0];
  assign s_496 = s_497 & s_499;
  assign s_497 = ~s_498;
  assign s_498 = s_489[1];
  assign s_499 = s_489[0];
  assign s_500 = s_501[1];
  assign s_501 = {s_502,s_508};
  assign s_502 = s_503 & s_506;
  assign s_503 = ~s_504;
  assign s_504 = s_505[1];
  assign s_505 = s_490[1:0];
  assign s_506 = ~s_507;
  assign s_507 = s_505[0];
  assign s_508 = s_509 & s_511;
  assign s_509 = ~s_510;
  assign s_510 = s_505[1];
  assign s_511 = s_505[0];
  assign s_512 = {s_513,s_515};
  assign s_513 = s_484 & s_514;
  assign s_514 = ~s_500;
  assign s_515 = s_484?s_516:s_517;
  assign s_516 = s_501[0:0];
  assign s_517 = s_485[0:0];
  assign s_518 = s_519[2];
  assign s_519 = {s_520,s_546};
  assign s_520 = s_521 & s_534;
  assign s_521 = s_522[1];
  assign s_522 = {s_523,s_530};
  assign s_523 = s_524 & s_528;
  assign s_524 = ~s_525;
  assign s_525 = s_526[1];
  assign s_526 = s_527[3:2];
  assign s_527 = s_491[3:0];
  assign s_528 = ~s_529;
  assign s_529 = s_526[0];
  assign s_530 = s_531 & s_533;
  assign s_531 = ~s_532;
  assign s_532 = s_526[1];
  assign s_533 = s_526[0];
  assign s_534 = s_535[1];
  assign s_535 = {s_536,s_542};
  assign s_536 = s_537 & s_540;
  assign s_537 = ~s_538;
  assign s_538 = s_539[1];
  assign s_539 = s_527[1:0];
  assign s_540 = ~s_541;
  assign s_541 = s_539[0];
  assign s_542 = s_543 & s_545;
  assign s_543 = ~s_544;
  assign s_544 = s_539[1];
  assign s_545 = s_539[0];
  assign s_546 = {s_547,s_549};
  assign s_547 = s_521 & s_548;
  assign s_548 = ~s_534;
  assign s_549 = s_521?s_550:s_551;
  assign s_550 = s_535[0:0];
  assign s_551 = s_522[0:0];
  assign s_552 = {s_553,s_555};
  assign s_553 = s_481 & s_554;
  assign s_554 = ~s_518;
  assign s_555 = s_481?s_556:s_557;
  assign s_556 = s_519[1:0];
  assign s_557 = s_482[1:0];
  assign s_558 = s_559[3];
  assign s_559 = {s_560,s_630};
  assign s_560 = s_561 & s_596;
  assign s_561 = s_562[2];
  assign s_562 = {s_563,s_590};
  assign s_563 = s_564 & s_578;
  assign s_564 = s_565[1];
  assign s_565 = {s_566,s_574};
  assign s_566 = s_567 & s_572;
  assign s_567 = ~s_568;
  assign s_568 = s_569[1];
  assign s_569 = s_570[3:2];
  assign s_570 = s_571[7:4];
  assign s_571 = s_492[7:0];
  assign s_572 = ~s_573;
  assign s_573 = s_569[0];
  assign s_574 = s_575 & s_577;
  assign s_575 = ~s_576;
  assign s_576 = s_569[1];
  assign s_577 = s_569[0];
  assign s_578 = s_579[1];
  assign s_579 = {s_580,s_586};
  assign s_580 = s_581 & s_584;
  assign s_581 = ~s_582;
  assign s_582 = s_583[1];
  assign s_583 = s_570[1:0];
  assign s_584 = ~s_585;
  assign s_585 = s_583[0];
  assign s_586 = s_587 & s_589;
  assign s_587 = ~s_588;
  assign s_588 = s_583[1];
  assign s_589 = s_583[0];
  assign s_590 = {s_591,s_593};
  assign s_591 = s_564 & s_592;
  assign s_592 = ~s_578;
  assign s_593 = s_564?s_594:s_595;
  assign s_594 = s_579[0:0];
  assign s_595 = s_565[0:0];
  assign s_596 = s_597[2];
  assign s_597 = {s_598,s_624};
  assign s_598 = s_599 & s_612;
  assign s_599 = s_600[1];
  assign s_600 = {s_601,s_608};
  assign s_601 = s_602 & s_606;
  assign s_602 = ~s_603;
  assign s_603 = s_604[1];
  assign s_604 = s_605[3:2];
  assign s_605 = s_571[3:0];
  assign s_606 = ~s_607;
  assign s_607 = s_604[0];
  assign s_608 = s_609 & s_611;
  assign s_609 = ~s_610;
  assign s_610 = s_604[1];
  assign s_611 = s_604[0];
  assign s_612 = s_613[1];
  assign s_613 = {s_614,s_620};
  assign s_614 = s_615 & s_618;
  assign s_615 = ~s_616;
  assign s_616 = s_617[1];
  assign s_617 = s_605[1:0];
  assign s_618 = ~s_619;
  assign s_619 = s_617[0];
  assign s_620 = s_621 & s_623;
  assign s_621 = ~s_622;
  assign s_622 = s_617[1];
  assign s_623 = s_617[0];
  assign s_624 = {s_625,s_627};
  assign s_625 = s_599 & s_626;
  assign s_626 = ~s_612;
  assign s_627 = s_599?s_628:s_629;
  assign s_628 = s_613[0:0];
  assign s_629 = s_600[0:0];
  assign s_630 = {s_631,s_633};
  assign s_631 = s_561 & s_632;
  assign s_632 = ~s_596;
  assign s_633 = s_561?s_634:s_635;
  assign s_634 = s_597[1:0];
  assign s_635 = s_562[1:0];
  assign s_636 = {s_637,s_639};
  assign s_637 = s_478 & s_638;
  assign s_638 = ~s_558;
  assign s_639 = s_478?s_640:s_641;
  assign s_640 = s_559[2:0];
  assign s_641 = s_479[2:0];
  assign s_642 = s_643[4];
  assign s_643 = {s_644,s_802};
  assign s_644 = s_645 & s_724;
  assign s_645 = s_646[3];
  assign s_646 = {s_647,s_718};
  assign s_647 = s_648 & s_684;
  assign s_648 = s_649[2];
  assign s_649 = {s_650,s_678};
  assign s_650 = s_651 & s_666;
  assign s_651 = s_652[1];
  assign s_652 = {s_653,s_662};
  assign s_653 = s_654 & s_660;
  assign s_654 = ~s_655;
  assign s_655 = s_656[1];
  assign s_656 = s_657[3:2];
  assign s_657 = s_658[7:4];
  assign s_658 = s_659[15:8];
  assign s_659 = s_493[15:0];
  assign s_660 = ~s_661;
  assign s_661 = s_656[0];
  assign s_662 = s_663 & s_665;
  assign s_663 = ~s_664;
  assign s_664 = s_656[1];
  assign s_665 = s_656[0];
  assign s_666 = s_667[1];
  assign s_667 = {s_668,s_674};
  assign s_668 = s_669 & s_672;
  assign s_669 = ~s_670;
  assign s_670 = s_671[1];
  assign s_671 = s_657[1:0];
  assign s_672 = ~s_673;
  assign s_673 = s_671[0];
  assign s_674 = s_675 & s_677;
  assign s_675 = ~s_676;
  assign s_676 = s_671[1];
  assign s_677 = s_671[0];
  assign s_678 = {s_679,s_681};
  assign s_679 = s_651 & s_680;
  assign s_680 = ~s_666;
  assign s_681 = s_651?s_682:s_683;
  assign s_682 = s_667[0:0];
  assign s_683 = s_652[0:0];
  assign s_684 = s_685[2];
  assign s_685 = {s_686,s_712};
  assign s_686 = s_687 & s_700;
  assign s_687 = s_688[1];
  assign s_688 = {s_689,s_696};
  assign s_689 = s_690 & s_694;
  assign s_690 = ~s_691;
  assign s_691 = s_692[1];
  assign s_692 = s_693[3:2];
  assign s_693 = s_658[3:0];
  assign s_694 = ~s_695;
  assign s_695 = s_692[0];
  assign s_696 = s_697 & s_699;
  assign s_697 = ~s_698;
  assign s_698 = s_692[1];
  assign s_699 = s_692[0];
  assign s_700 = s_701[1];
  assign s_701 = {s_702,s_708};
  assign s_702 = s_703 & s_706;
  assign s_703 = ~s_704;
  assign s_704 = s_705[1];
  assign s_705 = s_693[1:0];
  assign s_706 = ~s_707;
  assign s_707 = s_705[0];
  assign s_708 = s_709 & s_711;
  assign s_709 = ~s_710;
  assign s_710 = s_705[1];
  assign s_711 = s_705[0];
  assign s_712 = {s_713,s_715};
  assign s_713 = s_687 & s_714;
  assign s_714 = ~s_700;
  assign s_715 = s_687?s_716:s_717;
  assign s_716 = s_701[0:0];
  assign s_717 = s_688[0:0];
  assign s_718 = {s_719,s_721};
  assign s_719 = s_648 & s_720;
  assign s_720 = ~s_684;
  assign s_721 = s_648?s_722:s_723;
  assign s_722 = s_685[1:0];
  assign s_723 = s_649[1:0];
  assign s_724 = s_725[3];
  assign s_725 = {s_726,s_796};
  assign s_726 = s_727 & s_762;
  assign s_727 = s_728[2];
  assign s_728 = {s_729,s_756};
  assign s_729 = s_730 & s_744;
  assign s_730 = s_731[1];
  assign s_731 = {s_732,s_740};
  assign s_732 = s_733 & s_738;
  assign s_733 = ~s_734;
  assign s_734 = s_735[1];
  assign s_735 = s_736[3:2];
  assign s_736 = s_737[7:4];
  assign s_737 = s_659[7:0];
  assign s_738 = ~s_739;
  assign s_739 = s_735[0];
  assign s_740 = s_741 & s_743;
  assign s_741 = ~s_742;
  assign s_742 = s_735[1];
  assign s_743 = s_735[0];
  assign s_744 = s_745[1];
  assign s_745 = {s_746,s_752};
  assign s_746 = s_747 & s_750;
  assign s_747 = ~s_748;
  assign s_748 = s_749[1];
  assign s_749 = s_736[1:0];
  assign s_750 = ~s_751;
  assign s_751 = s_749[0];
  assign s_752 = s_753 & s_755;
  assign s_753 = ~s_754;
  assign s_754 = s_749[1];
  assign s_755 = s_749[0];
  assign s_756 = {s_757,s_759};
  assign s_757 = s_730 & s_758;
  assign s_758 = ~s_744;
  assign s_759 = s_730?s_760:s_761;
  assign s_760 = s_745[0:0];
  assign s_761 = s_731[0:0];
  assign s_762 = s_763[2];
  assign s_763 = {s_764,s_790};
  assign s_764 = s_765 & s_778;
  assign s_765 = s_766[1];
  assign s_766 = {s_767,s_774};
  assign s_767 = s_768 & s_772;
  assign s_768 = ~s_769;
  assign s_769 = s_770[1];
  assign s_770 = s_771[3:2];
  assign s_771 = s_737[3:0];
  assign s_772 = ~s_773;
  assign s_773 = s_770[0];
  assign s_774 = s_775 & s_777;
  assign s_775 = ~s_776;
  assign s_776 = s_770[1];
  assign s_777 = s_770[0];
  assign s_778 = s_779[1];
  assign s_779 = {s_780,s_786};
  assign s_780 = s_781 & s_784;
  assign s_781 = ~s_782;
  assign s_782 = s_783[1];
  assign s_783 = s_771[1:0];
  assign s_784 = ~s_785;
  assign s_785 = s_783[0];
  assign s_786 = s_787 & s_789;
  assign s_787 = ~s_788;
  assign s_788 = s_783[1];
  assign s_789 = s_783[0];
  assign s_790 = {s_791,s_793};
  assign s_791 = s_765 & s_792;
  assign s_792 = ~s_778;
  assign s_793 = s_765?s_794:s_795;
  assign s_794 = s_779[0:0];
  assign s_795 = s_766[0:0];
  assign s_796 = {s_797,s_799};
  assign s_797 = s_727 & s_798;
  assign s_798 = ~s_762;
  assign s_799 = s_727?s_800:s_801;
  assign s_800 = s_763[1:0];
  assign s_801 = s_728[1:0];
  assign s_802 = {s_803,s_805};
  assign s_803 = s_645 & s_804;
  assign s_804 = ~s_724;
  assign s_805 = s_645?s_806:s_807;
  assign s_806 = s_725[2:0];
  assign s_807 = s_646[2:0];
  assign s_808 = {s_809,s_811};
  assign s_809 = s_475 & s_810;
  assign s_810 = ~s_642;
  assign s_811 = s_475?s_812:s_813;
  assign s_812 = s_643[3:0];
  assign s_813 = s_476[3:0];
  assign s_814 = {s_815,s_817};
  assign s_815 = s_116 & s_816;
  assign s_816 = ~s_472;
  assign s_817 = s_116?s_818:s_819;
  assign s_818 = s_473[4:0];
  assign s_819 = s_117[4:0];
  dq #(12, 2) dq_s_820 (clk, s_820, s_821);
  assign s_821 = s_822 - s_827;
  dq #(12, 1) dq_s_822 (clk, s_822, s_823);
  assign s_823 = s_824 + s_826;
  assign s_824 = s_45?s_65:s_825;
  assign s_825 = s_66 + s_64;
  assign s_826 = 1'd1;
  assign s_827 = -12'd1022;
  assign s_828 = s_829 <= s_830;
  assign s_829 = s_113;
  dq #(12, 2) dq_s_830 (clk, s_830, s_821);
  assign s_831 = 1'd1;
  dq #(53, 1) dq_s_832 (clk, s_832, s_106);
  assign s_833 = s_834 & s_836;
  dq #(1, 1) dq_s_834 (clk, s_834, s_835);
  assign s_835 = s_107[3];
  assign s_836 = s_837 | s_844;
  assign s_837 = s_838 | s_840;
  dq #(1, 1) dq_s_838 (clk, s_838, s_839);
  assign s_839 = s_107[2];
  dq #(1, 1) dq_s_840 (clk, s_840, s_841);
  assign s_841 = s_842 | s_843;
  assign s_842 = s_107[1];
  assign s_843 = s_107[0];
  dq #(1, 1) dq_s_844 (clk, s_844, s_845);
  assign s_845 = s_106[0];
  assign s_846 = s_102[52:0];
  assign s_847 = s_102[53];
  assign s_848 = {s_849,s_860};
  assign s_849 = {s_850,s_851};
  dq #(1, 5) dq_s_850 (clk, s_850, s_3);
  assign s_851 = s_852 + s_859;
  assign s_852 = s_853[10:0];
  dq #(12, 1) dq_s_853 (clk, s_853, s_854);
  assign s_854 = s_855 + s_847;
  dq #(12, 1) dq_s_855 (clk, s_855, s_856);
  dq #(12, 1) dq_s_856 (clk, s_856, s_857);
  assign s_857 = s_858 - s_111;
  dq #(12, 3) dq_s_858 (clk, s_858, s_822);
  assign s_859 = 10'd1023;
  assign s_860 = s_99[51:0];
  assign s_861 = s_862 & s_864;
  assign s_862 = s_852 == s_863;
  assign s_863 = -11'd1022;
  assign s_864 = ~s_865;
  assign s_865 = s_99[52];
  assign s_866 = s_99 == s_867;
  assign s_867 = 53'd0;
  assign s_868 = s_869 | s_873;
  assign s_869 = s_870 | s_872;
  assign s_870 = $signed(s_853) > $signed(s_871);
  assign s_871 = 11'd1023;
  dq #(1, 7) dq_s_872 (clk, s_872, s_31);
  dq #(1, 7) dq_s_873 (clk, s_873, s_38);
  dq #(1, 7) dq_s_874 (clk, s_874, s_875);
  assign s_875 = s_876 | s_887;
  assign s_876 = s_877 | s_882;
  assign s_877 = s_878 & s_880;
  assign s_878 = s_18 == s_879;
  assign s_879 = 11'd1024;
  assign s_880 = s_35 != s_881;
  assign s_881 = 52'd0;
  assign s_882 = s_883 & s_885;
  assign s_883 = s_26 == s_884;
  assign s_884 = 11'd1024;
  assign s_885 = s_42 != s_886;
  assign s_886 = 52'd0;
  assign s_887 = s_31 & s_38;
  assign double_add_z = s_0;
endmodule
