module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module int_to_single(clk, int_to_single_a, int_to_single_z);
  input clk;
  input [31:0] int_to_single_a;
  output [31:0] int_to_single_z;
  wire [31:0] s_0;
  wire [31:0] s_1;
  wire [31:0] s_2;
  wire [0:0] s_3;
  wire [31:0] s_4;
  wire [30:0] s_5;
  wire [31:0] s_6;
  wire [31:0] s_7;
  wire [31:0] s_8;
  wire [30:0] s_9;
  wire [31:0] s_10;
  wire [31:0] s_11;
  wire [31:0] s_12;
  wire [30:0] s_13;
  wire [31:0] s_14;
  wire [31:0] s_15;
  wire [8:0] s_16;
  wire [8:0] s_17;
  wire [7:0] s_18;
  wire [22:0] s_19;
  wire [23:0] s_20;
  wire [23:0] s_21;
  wire [23:0] s_22;
  wire [24:0] s_23;
  wire [24:0] s_24;
  wire [24:0] s_25;
  wire [24:0] s_26;
  wire [23:0] s_27;
  wire [31:0] s_28;
  wire [31:0] s_29;
  wire [31:0] s_30;
  wire [31:0] s_31;
  wire [31:0] s_32;
  wire [31:0] s_33;
  wire [5:0] s_34;
  wire [5:0] s_35;
  wire [0:0] s_36;
  wire [0:0] s_37;
  wire [4:0] s_38;
  wire [0:0] s_39;
  wire [0:0] s_40;
  wire [3:0] s_41;
  wire [0:0] s_42;
  wire [0:0] s_43;
  wire [2:0] s_44;
  wire [0:0] s_45;
  wire [0:0] s_46;
  wire [1:0] s_47;
  wire [0:0] s_48;
  wire [0:0] s_49;
  wire [0:0] s_50;
  wire [1:0] s_51;
  wire [3:0] s_52;
  wire [7:0] s_53;
  wire [15:0] s_54;
  wire [0:0] s_55;
  wire [0:0] s_56;
  wire [0:0] s_57;
  wire [0:0] s_58;
  wire [0:0] s_59;
  wire [0:0] s_60;
  wire [0:0] s_61;
  wire [1:0] s_62;
  wire [0:0] s_63;
  wire [0:0] s_64;
  wire [0:0] s_65;
  wire [1:0] s_66;
  wire [0:0] s_67;
  wire [0:0] s_68;
  wire [0:0] s_69;
  wire [0:0] s_70;
  wire [0:0] s_71;
  wire [0:0] s_72;
  wire [1:0] s_73;
  wire [0:0] s_74;
  wire [0:0] s_75;
  wire [0:0] s_76;
  wire [0:0] s_77;
  wire [0:0] s_78;
  wire [0:0] s_79;
  wire [2:0] s_80;
  wire [0:0] s_81;
  wire [0:0] s_82;
  wire [1:0] s_83;
  wire [0:0] s_84;
  wire [0:0] s_85;
  wire [0:0] s_86;
  wire [1:0] s_87;
  wire [3:0] s_88;
  wire [0:0] s_89;
  wire [0:0] s_90;
  wire [0:0] s_91;
  wire [0:0] s_92;
  wire [0:0] s_93;
  wire [0:0] s_94;
  wire [0:0] s_95;
  wire [1:0] s_96;
  wire [0:0] s_97;
  wire [0:0] s_98;
  wire [0:0] s_99;
  wire [1:0] s_100;
  wire [0:0] s_101;
  wire [0:0] s_102;
  wire [0:0] s_103;
  wire [0:0] s_104;
  wire [0:0] s_105;
  wire [0:0] s_106;
  wire [1:0] s_107;
  wire [0:0] s_108;
  wire [0:0] s_109;
  wire [0:0] s_110;
  wire [0:0] s_111;
  wire [0:0] s_112;
  wire [2:0] s_113;
  wire [0:0] s_114;
  wire [0:0] s_115;
  wire [1:0] s_116;
  wire [1:0] s_117;
  wire [1:0] s_118;
  wire [0:0] s_119;
  wire [3:0] s_120;
  wire [0:0] s_121;
  wire [0:0] s_122;
  wire [2:0] s_123;
  wire [0:0] s_124;
  wire [0:0] s_125;
  wire [1:0] s_126;
  wire [0:0] s_127;
  wire [0:0] s_128;
  wire [0:0] s_129;
  wire [1:0] s_130;
  wire [3:0] s_131;
  wire [7:0] s_132;
  wire [0:0] s_133;
  wire [0:0] s_134;
  wire [0:0] s_135;
  wire [0:0] s_136;
  wire [0:0] s_137;
  wire [0:0] s_138;
  wire [0:0] s_139;
  wire [1:0] s_140;
  wire [0:0] s_141;
  wire [0:0] s_142;
  wire [0:0] s_143;
  wire [1:0] s_144;
  wire [0:0] s_145;
  wire [0:0] s_146;
  wire [0:0] s_147;
  wire [0:0] s_148;
  wire [0:0] s_149;
  wire [0:0] s_150;
  wire [1:0] s_151;
  wire [0:0] s_152;
  wire [0:0] s_153;
  wire [0:0] s_154;
  wire [0:0] s_155;
  wire [0:0] s_156;
  wire [0:0] s_157;
  wire [2:0] s_158;
  wire [0:0] s_159;
  wire [0:0] s_160;
  wire [1:0] s_161;
  wire [0:0] s_162;
  wire [0:0] s_163;
  wire [0:0] s_164;
  wire [1:0] s_165;
  wire [3:0] s_166;
  wire [0:0] s_167;
  wire [0:0] s_168;
  wire [0:0] s_169;
  wire [0:0] s_170;
  wire [0:0] s_171;
  wire [0:0] s_172;
  wire [0:0] s_173;
  wire [1:0] s_174;
  wire [0:0] s_175;
  wire [0:0] s_176;
  wire [0:0] s_177;
  wire [1:0] s_178;
  wire [0:0] s_179;
  wire [0:0] s_180;
  wire [0:0] s_181;
  wire [0:0] s_182;
  wire [0:0] s_183;
  wire [0:0] s_184;
  wire [1:0] s_185;
  wire [0:0] s_186;
  wire [0:0] s_187;
  wire [0:0] s_188;
  wire [0:0] s_189;
  wire [0:0] s_190;
  wire [2:0] s_191;
  wire [0:0] s_192;
  wire [0:0] s_193;
  wire [1:0] s_194;
  wire [1:0] s_195;
  wire [1:0] s_196;
  wire [3:0] s_197;
  wire [0:0] s_198;
  wire [0:0] s_199;
  wire [2:0] s_200;
  wire [2:0] s_201;
  wire [2:0] s_202;
  wire [0:0] s_203;
  wire [4:0] s_204;
  wire [0:0] s_205;
  wire [0:0] s_206;
  wire [3:0] s_207;
  wire [0:0] s_208;
  wire [0:0] s_209;
  wire [2:0] s_210;
  wire [0:0] s_211;
  wire [0:0] s_212;
  wire [1:0] s_213;
  wire [0:0] s_214;
  wire [0:0] s_215;
  wire [0:0] s_216;
  wire [1:0] s_217;
  wire [3:0] s_218;
  wire [7:0] s_219;
  wire [15:0] s_220;
  wire [0:0] s_221;
  wire [0:0] s_222;
  wire [0:0] s_223;
  wire [0:0] s_224;
  wire [0:0] s_225;
  wire [0:0] s_226;
  wire [0:0] s_227;
  wire [1:0] s_228;
  wire [0:0] s_229;
  wire [0:0] s_230;
  wire [0:0] s_231;
  wire [1:0] s_232;
  wire [0:0] s_233;
  wire [0:0] s_234;
  wire [0:0] s_235;
  wire [0:0] s_236;
  wire [0:0] s_237;
  wire [0:0] s_238;
  wire [1:0] s_239;
  wire [0:0] s_240;
  wire [0:0] s_241;
  wire [0:0] s_242;
  wire [0:0] s_243;
  wire [0:0] s_244;
  wire [0:0] s_245;
  wire [2:0] s_246;
  wire [0:0] s_247;
  wire [0:0] s_248;
  wire [1:0] s_249;
  wire [0:0] s_250;
  wire [0:0] s_251;
  wire [0:0] s_252;
  wire [1:0] s_253;
  wire [3:0] s_254;
  wire [0:0] s_255;
  wire [0:0] s_256;
  wire [0:0] s_257;
  wire [0:0] s_258;
  wire [0:0] s_259;
  wire [0:0] s_260;
  wire [0:0] s_261;
  wire [1:0] s_262;
  wire [0:0] s_263;
  wire [0:0] s_264;
  wire [0:0] s_265;
  wire [1:0] s_266;
  wire [0:0] s_267;
  wire [0:0] s_268;
  wire [0:0] s_269;
  wire [0:0] s_270;
  wire [0:0] s_271;
  wire [0:0] s_272;
  wire [1:0] s_273;
  wire [0:0] s_274;
  wire [0:0] s_275;
  wire [0:0] s_276;
  wire [0:0] s_277;
  wire [0:0] s_278;
  wire [2:0] s_279;
  wire [0:0] s_280;
  wire [0:0] s_281;
  wire [1:0] s_282;
  wire [1:0] s_283;
  wire [1:0] s_284;
  wire [0:0] s_285;
  wire [3:0] s_286;
  wire [0:0] s_287;
  wire [0:0] s_288;
  wire [2:0] s_289;
  wire [0:0] s_290;
  wire [0:0] s_291;
  wire [1:0] s_292;
  wire [0:0] s_293;
  wire [0:0] s_294;
  wire [0:0] s_295;
  wire [1:0] s_296;
  wire [3:0] s_297;
  wire [7:0] s_298;
  wire [0:0] s_299;
  wire [0:0] s_300;
  wire [0:0] s_301;
  wire [0:0] s_302;
  wire [0:0] s_303;
  wire [0:0] s_304;
  wire [0:0] s_305;
  wire [1:0] s_306;
  wire [0:0] s_307;
  wire [0:0] s_308;
  wire [0:0] s_309;
  wire [1:0] s_310;
  wire [0:0] s_311;
  wire [0:0] s_312;
  wire [0:0] s_313;
  wire [0:0] s_314;
  wire [0:0] s_315;
  wire [0:0] s_316;
  wire [1:0] s_317;
  wire [0:0] s_318;
  wire [0:0] s_319;
  wire [0:0] s_320;
  wire [0:0] s_321;
  wire [0:0] s_322;
  wire [0:0] s_323;
  wire [2:0] s_324;
  wire [0:0] s_325;
  wire [0:0] s_326;
  wire [1:0] s_327;
  wire [0:0] s_328;
  wire [0:0] s_329;
  wire [0:0] s_330;
  wire [1:0] s_331;
  wire [3:0] s_332;
  wire [0:0] s_333;
  wire [0:0] s_334;
  wire [0:0] s_335;
  wire [0:0] s_336;
  wire [0:0] s_337;
  wire [0:0] s_338;
  wire [0:0] s_339;
  wire [1:0] s_340;
  wire [0:0] s_341;
  wire [0:0] s_342;
  wire [0:0] s_343;
  wire [1:0] s_344;
  wire [0:0] s_345;
  wire [0:0] s_346;
  wire [0:0] s_347;
  wire [0:0] s_348;
  wire [0:0] s_349;
  wire [0:0] s_350;
  wire [1:0] s_351;
  wire [0:0] s_352;
  wire [0:0] s_353;
  wire [0:0] s_354;
  wire [0:0] s_355;
  wire [0:0] s_356;
  wire [2:0] s_357;
  wire [0:0] s_358;
  wire [0:0] s_359;
  wire [1:0] s_360;
  wire [1:0] s_361;
  wire [1:0] s_362;
  wire [3:0] s_363;
  wire [0:0] s_364;
  wire [0:0] s_365;
  wire [2:0] s_366;
  wire [2:0] s_367;
  wire [2:0] s_368;
  wire [4:0] s_369;
  wire [0:0] s_370;
  wire [0:0] s_371;
  wire [3:0] s_372;
  wire [3:0] s_373;
  wire [3:0] s_374;
  wire [0:0] s_375;
  wire [23:0] s_376;
  wire [0:0] s_377;
  wire [0:0] s_378;
  wire [0:0] s_379;
  wire [0:0] s_380;
  wire [0:0] s_381;
  wire [0:0] s_382;
  wire [0:0] s_383;
  wire [0:0] s_384;
  wire [0:0] s_385;
  wire [5:0] s_386;
  wire [0:0] s_387;
  wire [0:0] s_388;
  wire [0:0] s_389;
  wire [23:0] s_390;
  wire [0:0] s_391;
  wire [31:0] s_392;
  wire [8:0] s_393;
  wire [0:0] s_394;
  wire [7:0] s_395;
  wire [7:0] s_396;
  wire [7:0] s_397;
  wire [7:0] s_398;
  wire [7:0] s_399;
  wire [7:0] s_400;
  wire [6:0] s_401;
  wire [22:0] s_402;
  wire [0:0] s_403;
  wire [0:0] s_404;
  wire [7:0] s_405;
  wire [0:0] s_406;
  wire [0:0] s_407;
  wire [0:0] s_408;
  wire [23:0] s_409;
  wire [0:0] s_410;
  wire [0:0] s_411;

  assign s_0 = s_411?s_1:s_6;
  dq #(32, 5) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_5};
  assign s_3 = s_4[31];
  assign s_4 = int_to_single_a;
  assign s_5 = 31'd2143289344;
  assign s_6 = s_410?s_7:s_10;
  dq #(32, 5) dq_s_7 (clk, s_7, s_8);
  assign s_8 = {s_3,s_9};
  assign s_9 = 31'd2139095040;
  assign s_10 = s_408?s_11:s_14;
  dq #(32, 5) dq_s_11 (clk, s_11, s_12);
  assign s_12 = {s_3,s_13};
  assign s_13 = 31'd0;
  assign s_14 = s_403?s_15:s_392;
  assign s_15 = {s_16,s_19};
  dq #(9, 5) dq_s_16 (clk, s_16, s_17);
  assign s_17 = {s_3,s_18};
  assign s_18 = 8'd0;
  assign s_19 = s_20[22:0];
  dq #(24, 1) dq_s_20 (clk, s_20, s_21);
  assign s_21 = s_391?s_22:s_390;
  assign s_22 = s_23[24:1];
  assign s_23 = s_377?s_24:s_376;
  dq #(25, 1) dq_s_24 (clk, s_24, s_25);
  assign s_25 = s_26 + s_375;
  assign s_26 = s_27;
  assign s_27 = s_28[31:8];
  dq #(32, 1) dq_s_28 (clk, s_28, s_29);
  assign s_29 = s_30 << s_34;
  dq #(32, 1) dq_s_30 (clk, s_30, s_31);
  dq #(32, 1) dq_s_31 (clk, s_31, s_32);
  assign s_32 = s_3?s_33:s_4;
  assign s_33 = -s_4;
  dq #(6, 1) dq_s_34 (clk, s_34, s_35);
  assign s_35 = {s_36,s_369};
  assign s_36 = s_37 & s_203;
  assign s_37 = s_38[4];
  assign s_38 = {s_39,s_197};
  assign s_39 = s_40 & s_119;
  assign s_40 = s_41[3];
  assign s_41 = {s_42,s_113};
  assign s_42 = s_43 & s_79;
  assign s_43 = s_44[2];
  assign s_44 = {s_45,s_73};
  assign s_45 = s_46 & s_61;
  assign s_46 = s_47[1];
  assign s_47 = {s_48,s_57};
  assign s_48 = s_49 & s_55;
  assign s_49 = ~s_50;
  assign s_50 = s_51[1];
  assign s_51 = s_52[3:2];
  assign s_52 = s_53[7:4];
  assign s_53 = s_54[15:8];
  assign s_54 = s_31[31:16];
  assign s_55 = ~s_56;
  assign s_56 = s_51[0];
  assign s_57 = s_58 & s_60;
  assign s_58 = ~s_59;
  assign s_59 = s_51[1];
  assign s_60 = s_51[0];
  assign s_61 = s_62[1];
  assign s_62 = {s_63,s_69};
  assign s_63 = s_64 & s_67;
  assign s_64 = ~s_65;
  assign s_65 = s_66[1];
  assign s_66 = s_52[1:0];
  assign s_67 = ~s_68;
  assign s_68 = s_66[0];
  assign s_69 = s_70 & s_72;
  assign s_70 = ~s_71;
  assign s_71 = s_66[1];
  assign s_72 = s_66[0];
  assign s_73 = {s_74,s_76};
  assign s_74 = s_46 & s_75;
  assign s_75 = ~s_61;
  assign s_76 = s_46?s_77:s_78;
  assign s_77 = s_62[0:0];
  assign s_78 = s_47[0:0];
  assign s_79 = s_80[2];
  assign s_80 = {s_81,s_107};
  assign s_81 = s_82 & s_95;
  assign s_82 = s_83[1];
  assign s_83 = {s_84,s_91};
  assign s_84 = s_85 & s_89;
  assign s_85 = ~s_86;
  assign s_86 = s_87[1];
  assign s_87 = s_88[3:2];
  assign s_88 = s_53[3:0];
  assign s_89 = ~s_90;
  assign s_90 = s_87[0];
  assign s_91 = s_92 & s_94;
  assign s_92 = ~s_93;
  assign s_93 = s_87[1];
  assign s_94 = s_87[0];
  assign s_95 = s_96[1];
  assign s_96 = {s_97,s_103};
  assign s_97 = s_98 & s_101;
  assign s_98 = ~s_99;
  assign s_99 = s_100[1];
  assign s_100 = s_88[1:0];
  assign s_101 = ~s_102;
  assign s_102 = s_100[0];
  assign s_103 = s_104 & s_106;
  assign s_104 = ~s_105;
  assign s_105 = s_100[1];
  assign s_106 = s_100[0];
  assign s_107 = {s_108,s_110};
  assign s_108 = s_82 & s_109;
  assign s_109 = ~s_95;
  assign s_110 = s_82?s_111:s_112;
  assign s_111 = s_96[0:0];
  assign s_112 = s_83[0:0];
  assign s_113 = {s_114,s_116};
  assign s_114 = s_43 & s_115;
  assign s_115 = ~s_79;
  assign s_116 = s_43?s_117:s_118;
  assign s_117 = s_80[1:0];
  assign s_118 = s_44[1:0];
  assign s_119 = s_120[3];
  assign s_120 = {s_121,s_191};
  assign s_121 = s_122 & s_157;
  assign s_122 = s_123[2];
  assign s_123 = {s_124,s_151};
  assign s_124 = s_125 & s_139;
  assign s_125 = s_126[1];
  assign s_126 = {s_127,s_135};
  assign s_127 = s_128 & s_133;
  assign s_128 = ~s_129;
  assign s_129 = s_130[1];
  assign s_130 = s_131[3:2];
  assign s_131 = s_132[7:4];
  assign s_132 = s_54[7:0];
  assign s_133 = ~s_134;
  assign s_134 = s_130[0];
  assign s_135 = s_136 & s_138;
  assign s_136 = ~s_137;
  assign s_137 = s_130[1];
  assign s_138 = s_130[0];
  assign s_139 = s_140[1];
  assign s_140 = {s_141,s_147};
  assign s_141 = s_142 & s_145;
  assign s_142 = ~s_143;
  assign s_143 = s_144[1];
  assign s_144 = s_131[1:0];
  assign s_145 = ~s_146;
  assign s_146 = s_144[0];
  assign s_147 = s_148 & s_150;
  assign s_148 = ~s_149;
  assign s_149 = s_144[1];
  assign s_150 = s_144[0];
  assign s_151 = {s_152,s_154};
  assign s_152 = s_125 & s_153;
  assign s_153 = ~s_139;
  assign s_154 = s_125?s_155:s_156;
  assign s_155 = s_140[0:0];
  assign s_156 = s_126[0:0];
  assign s_157 = s_158[2];
  assign s_158 = {s_159,s_185};
  assign s_159 = s_160 & s_173;
  assign s_160 = s_161[1];
  assign s_161 = {s_162,s_169};
  assign s_162 = s_163 & s_167;
  assign s_163 = ~s_164;
  assign s_164 = s_165[1];
  assign s_165 = s_166[3:2];
  assign s_166 = s_132[3:0];
  assign s_167 = ~s_168;
  assign s_168 = s_165[0];
  assign s_169 = s_170 & s_172;
  assign s_170 = ~s_171;
  assign s_171 = s_165[1];
  assign s_172 = s_165[0];
  assign s_173 = s_174[1];
  assign s_174 = {s_175,s_181};
  assign s_175 = s_176 & s_179;
  assign s_176 = ~s_177;
  assign s_177 = s_178[1];
  assign s_178 = s_166[1:0];
  assign s_179 = ~s_180;
  assign s_180 = s_178[0];
  assign s_181 = s_182 & s_184;
  assign s_182 = ~s_183;
  assign s_183 = s_178[1];
  assign s_184 = s_178[0];
  assign s_185 = {s_186,s_188};
  assign s_186 = s_160 & s_187;
  assign s_187 = ~s_173;
  assign s_188 = s_160?s_189:s_190;
  assign s_189 = s_174[0:0];
  assign s_190 = s_161[0:0];
  assign s_191 = {s_192,s_194};
  assign s_192 = s_122 & s_193;
  assign s_193 = ~s_157;
  assign s_194 = s_122?s_195:s_196;
  assign s_195 = s_158[1:0];
  assign s_196 = s_123[1:0];
  assign s_197 = {s_198,s_200};
  assign s_198 = s_40 & s_199;
  assign s_199 = ~s_119;
  assign s_200 = s_40?s_201:s_202;
  assign s_201 = s_120[2:0];
  assign s_202 = s_41[2:0];
  assign s_203 = s_204[4];
  assign s_204 = {s_205,s_363};
  assign s_205 = s_206 & s_285;
  assign s_206 = s_207[3];
  assign s_207 = {s_208,s_279};
  assign s_208 = s_209 & s_245;
  assign s_209 = s_210[2];
  assign s_210 = {s_211,s_239};
  assign s_211 = s_212 & s_227;
  assign s_212 = s_213[1];
  assign s_213 = {s_214,s_223};
  assign s_214 = s_215 & s_221;
  assign s_215 = ~s_216;
  assign s_216 = s_217[1];
  assign s_217 = s_218[3:2];
  assign s_218 = s_219[7:4];
  assign s_219 = s_220[15:8];
  assign s_220 = s_31[15:0];
  assign s_221 = ~s_222;
  assign s_222 = s_217[0];
  assign s_223 = s_224 & s_226;
  assign s_224 = ~s_225;
  assign s_225 = s_217[1];
  assign s_226 = s_217[0];
  assign s_227 = s_228[1];
  assign s_228 = {s_229,s_235};
  assign s_229 = s_230 & s_233;
  assign s_230 = ~s_231;
  assign s_231 = s_232[1];
  assign s_232 = s_218[1:0];
  assign s_233 = ~s_234;
  assign s_234 = s_232[0];
  assign s_235 = s_236 & s_238;
  assign s_236 = ~s_237;
  assign s_237 = s_232[1];
  assign s_238 = s_232[0];
  assign s_239 = {s_240,s_242};
  assign s_240 = s_212 & s_241;
  assign s_241 = ~s_227;
  assign s_242 = s_212?s_243:s_244;
  assign s_243 = s_228[0:0];
  assign s_244 = s_213[0:0];
  assign s_245 = s_246[2];
  assign s_246 = {s_247,s_273};
  assign s_247 = s_248 & s_261;
  assign s_248 = s_249[1];
  assign s_249 = {s_250,s_257};
  assign s_250 = s_251 & s_255;
  assign s_251 = ~s_252;
  assign s_252 = s_253[1];
  assign s_253 = s_254[3:2];
  assign s_254 = s_219[3:0];
  assign s_255 = ~s_256;
  assign s_256 = s_253[0];
  assign s_257 = s_258 & s_260;
  assign s_258 = ~s_259;
  assign s_259 = s_253[1];
  assign s_260 = s_253[0];
  assign s_261 = s_262[1];
  assign s_262 = {s_263,s_269};
  assign s_263 = s_264 & s_267;
  assign s_264 = ~s_265;
  assign s_265 = s_266[1];
  assign s_266 = s_254[1:0];
  assign s_267 = ~s_268;
  assign s_268 = s_266[0];
  assign s_269 = s_270 & s_272;
  assign s_270 = ~s_271;
  assign s_271 = s_266[1];
  assign s_272 = s_266[0];
  assign s_273 = {s_274,s_276};
  assign s_274 = s_248 & s_275;
  assign s_275 = ~s_261;
  assign s_276 = s_248?s_277:s_278;
  assign s_277 = s_262[0:0];
  assign s_278 = s_249[0:0];
  assign s_279 = {s_280,s_282};
  assign s_280 = s_209 & s_281;
  assign s_281 = ~s_245;
  assign s_282 = s_209?s_283:s_284;
  assign s_283 = s_246[1:0];
  assign s_284 = s_210[1:0];
  assign s_285 = s_286[3];
  assign s_286 = {s_287,s_357};
  assign s_287 = s_288 & s_323;
  assign s_288 = s_289[2];
  assign s_289 = {s_290,s_317};
  assign s_290 = s_291 & s_305;
  assign s_291 = s_292[1];
  assign s_292 = {s_293,s_301};
  assign s_293 = s_294 & s_299;
  assign s_294 = ~s_295;
  assign s_295 = s_296[1];
  assign s_296 = s_297[3:2];
  assign s_297 = s_298[7:4];
  assign s_298 = s_220[7:0];
  assign s_299 = ~s_300;
  assign s_300 = s_296[0];
  assign s_301 = s_302 & s_304;
  assign s_302 = ~s_303;
  assign s_303 = s_296[1];
  assign s_304 = s_296[0];
  assign s_305 = s_306[1];
  assign s_306 = {s_307,s_313};
  assign s_307 = s_308 & s_311;
  assign s_308 = ~s_309;
  assign s_309 = s_310[1];
  assign s_310 = s_297[1:0];
  assign s_311 = ~s_312;
  assign s_312 = s_310[0];
  assign s_313 = s_314 & s_316;
  assign s_314 = ~s_315;
  assign s_315 = s_310[1];
  assign s_316 = s_310[0];
  assign s_317 = {s_318,s_320};
  assign s_318 = s_291 & s_319;
  assign s_319 = ~s_305;
  assign s_320 = s_291?s_321:s_322;
  assign s_321 = s_306[0:0];
  assign s_322 = s_292[0:0];
  assign s_323 = s_324[2];
  assign s_324 = {s_325,s_351};
  assign s_325 = s_326 & s_339;
  assign s_326 = s_327[1];
  assign s_327 = {s_328,s_335};
  assign s_328 = s_329 & s_333;
  assign s_329 = ~s_330;
  assign s_330 = s_331[1];
  assign s_331 = s_332[3:2];
  assign s_332 = s_298[3:0];
  assign s_333 = ~s_334;
  assign s_334 = s_331[0];
  assign s_335 = s_336 & s_338;
  assign s_336 = ~s_337;
  assign s_337 = s_331[1];
  assign s_338 = s_331[0];
  assign s_339 = s_340[1];
  assign s_340 = {s_341,s_347};
  assign s_341 = s_342 & s_345;
  assign s_342 = ~s_343;
  assign s_343 = s_344[1];
  assign s_344 = s_332[1:0];
  assign s_345 = ~s_346;
  assign s_346 = s_344[0];
  assign s_347 = s_348 & s_350;
  assign s_348 = ~s_349;
  assign s_349 = s_344[1];
  assign s_350 = s_344[0];
  assign s_351 = {s_352,s_354};
  assign s_352 = s_326 & s_353;
  assign s_353 = ~s_339;
  assign s_354 = s_326?s_355:s_356;
  assign s_355 = s_340[0:0];
  assign s_356 = s_327[0:0];
  assign s_357 = {s_358,s_360};
  assign s_358 = s_288 & s_359;
  assign s_359 = ~s_323;
  assign s_360 = s_288?s_361:s_362;
  assign s_361 = s_324[1:0];
  assign s_362 = s_289[1:0];
  assign s_363 = {s_364,s_366};
  assign s_364 = s_206 & s_365;
  assign s_365 = ~s_285;
  assign s_366 = s_206?s_367:s_368;
  assign s_367 = s_286[2:0];
  assign s_368 = s_207[2:0];
  assign s_369 = {s_370,s_372};
  assign s_370 = s_37 & s_371;
  assign s_371 = ~s_203;
  assign s_372 = s_37?s_373:s_374;
  assign s_373 = s_204[3:0];
  assign s_374 = s_38[3:0];
  assign s_375 = 1'd1;
  dq #(24, 1) dq_s_376 (clk, s_376, s_27);
  assign s_377 = s_378 & s_380;
  dq #(1, 1) dq_s_378 (clk, s_378, s_379);
  assign s_379 = s_28[7];
  assign s_380 = s_381 | s_388;
  assign s_381 = s_382 | s_384;
  dq #(1, 1) dq_s_382 (clk, s_382, s_383);
  assign s_383 = s_28[6];
  dq #(1, 1) dq_s_384 (clk, s_384, s_385);
  assign s_385 = s_386 != s_387;
  assign s_386 = s_28[5:0];
  assign s_387 = 1'd0;
  dq #(1, 1) dq_s_388 (clk, s_388, s_389);
  assign s_389 = s_27[0];
  assign s_390 = s_23[23:0];
  assign s_391 = s_23[24];
  assign s_392 = {s_393,s_402};
  assign s_393 = {s_394,s_395};
  dq #(1, 5) dq_s_394 (clk, s_394, s_3);
  assign s_395 = s_396 + s_401;
  dq #(8, 1) dq_s_396 (clk, s_396, s_397);
  assign s_397 = s_398 + s_391;
  dq #(8, 2) dq_s_398 (clk, s_398, s_399);
  assign s_399 = s_400 - s_34;
  assign s_400 = 8'd31;
  assign s_401 = 7'd127;
  assign s_402 = s_20[22:0];
  assign s_403 = s_404 & s_406;
  assign s_404 = s_396 == s_405;
  assign s_405 = -8'd126;
  assign s_406 = ~s_407;
  assign s_407 = s_20[23];
  assign s_408 = s_20 == s_409;
  assign s_409 = 24'd0;
  assign s_410 = 1'd0;
  assign s_411 = 1'd0;
  assign int_to_single_z = s_0;
endmodule
