module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module double_mul(clk, double_mul_a, double_mul_b, double_mul_z);
  input clk;
  input [63:0] double_mul_a;
  input [63:0] double_mul_b;
  output [63:0] double_mul_z;
  wire [63:0] s_0;
  wire [63:0] s_1;
  wire [63:0] s_2;
  wire [0:0] s_3;
  wire [0:0] s_4;
  wire [63:0] s_5;
  wire [0:0] s_6;
  wire [63:0] s_7;
  wire [62:0] s_8;
  wire [63:0] s_9;
  wire [63:0] s_10;
  wire [63:0] s_11;
  wire [62:0] s_12;
  wire [63:0] s_13;
  wire [63:0] s_14;
  wire [63:0] s_15;
  wire [62:0] s_16;
  wire [63:0] s_17;
  wire [63:0] s_18;
  wire [11:0] s_19;
  wire [11:0] s_20;
  wire [10:0] s_21;
  wire [51:0] s_22;
  wire [52:0] s_23;
  wire [52:0] s_24;
  wire [52:0] s_25;
  wire [53:0] s_26;
  wire [53:0] s_27;
  wire [53:0] s_28;
  wire [53:0] s_29;
  wire [52:0] s_30;
  wire [105:0] s_31;
  wire [105:0] s_32;
  wire [105:0] s_33;
  wire [105:0] s_34;
  wire [105:0] s_35;
  wire [105:0] s_36;
  wire [118:0] s_37;
  wire [16:0] s_38;
  wire [48:0] s_39;
  wire [48:0] s_40;
  wire [47:0] s_41;
  wire [33:0] s_42;
  wire [33:0] s_43;
  wire [33:0] s_44;
  wire [16:0] s_45;
  wire [67:0] s_46;
  wire [52:0] s_47;
  wire [0:0] s_48;
  wire [0:0] s_49;
  wire [0:0] s_50;
  wire [0:0] s_51;
  wire [10:0] s_52;
  wire [10:0] s_53;
  wire [9:0] s_54;
  wire [10:0] s_55;
  wire [51:0] s_56;
  wire [16:0] s_57;
  wire [67:0] s_58;
  wire [52:0] s_59;
  wire [0:0] s_60;
  wire [0:0] s_61;
  wire [0:0] s_62;
  wire [0:0] s_63;
  wire [10:0] s_64;
  wire [10:0] s_65;
  wire [9:0] s_66;
  wire [10:0] s_67;
  wire [51:0] s_68;
  wire [47:0] s_69;
  wire [47:0] s_70;
  wire [47:0] s_71;
  wire [46:0] s_72;
  wire [33:0] s_73;
  wire [33:0] s_74;
  wire [33:0] s_75;
  wire [16:0] s_76;
  wire [46:0] s_77;
  wire [46:0] s_78;
  wire [45:0] s_79;
  wire [33:0] s_80;
  wire [33:0] s_81;
  wire [33:0] s_82;
  wire [16:0] s_83;
  wire [45:0] s_84;
  wire [45:0] s_85;
  wire [45:0] s_86;
  wire [44:0] s_87;
  wire [33:0] s_88;
  wire [33:0] s_89;
  wire [33:0] s_90;
  wire [16:0] s_91;
  wire [44:0] s_92;
  wire [44:0] s_93;
  wire [43:0] s_94;
  wire [33:0] s_95;
  wire [33:0] s_96;
  wire [33:0] s_97;
  wire [43:0] s_98;
  wire [43:0] s_99;
  wire [42:0] s_100;
  wire [33:0] s_101;
  wire [33:0] s_102;
  wire [33:0] s_103;
  wire [16:0] s_104;
  wire [42:0] s_105;
  wire [42:0] s_106;
  wire [42:0] s_107;
  wire [41:0] s_108;
  wire [33:0] s_109;
  wire [33:0] s_110;
  wire [33:0] s_111;
  wire [16:0] s_112;
  wire [41:0] s_113;
  wire [41:0] s_114;
  wire [40:0] s_115;
  wire [33:0] s_116;
  wire [33:0] s_117;
  wire [33:0] s_118;
  wire [40:0] s_119;
  wire [40:0] s_120;
  wire [39:0] s_121;
  wire [33:0] s_122;
  wire [33:0] s_123;
  wire [33:0] s_124;
  wire [39:0] s_125;
  wire [39:0] s_126;
  wire [38:0] s_127;
  wire [33:0] s_128;
  wire [33:0] s_129;
  wire [33:0] s_130;
  wire [16:0] s_131;
  wire [38:0] s_132;
  wire [38:0] s_133;
  wire [38:0] s_134;
  wire [37:0] s_135;
  wire [33:0] s_136;
  wire [33:0] s_137;
  wire [33:0] s_138;
  wire [37:0] s_139;
  wire [37:0] s_140;
  wire [36:0] s_141;
  wire [33:0] s_142;
  wire [33:0] s_143;
  wire [33:0] s_144;
  wire [36:0] s_145;
  wire [36:0] s_146;
  wire [35:0] s_147;
  wire [33:0] s_148;
  wire [33:0] s_149;
  wire [33:0] s_150;
  wire [35:0] s_151;
  wire [35:0] s_152;
  wire [35:0] s_153;
  wire [34:0] s_154;
  wire [33:0] s_155;
  wire [33:0] s_156;
  wire [33:0] s_157;
  wire [34:0] s_158;
  wire [34:0] s_159;
  wire [33:0] s_160;
  wire [33:0] s_161;
  wire [33:0] s_162;
  wire [33:0] s_163;
  wire [33:0] s_164;
  wire [33:0] s_165;
  wire [4:0] s_166;
  wire [4:0] s_167;
  wire [4:0] s_168;
  wire [4:0] s_169;
  wire [4:0] s_170;
  wire [4:0] s_171;
  wire [101:0] s_172;
  wire [101:0] s_173;
  wire [16:0] s_174;
  wire [84:0] s_175;
  wire [84:0] s_176;
  wire [16:0] s_177;
  wire [67:0] s_178;
  wire [67:0] s_179;
  wire [16:0] s_180;
  wire [50:0] s_181;
  wire [50:0] s_182;
  wire [16:0] s_183;
  wire [33:0] s_184;
  wire [33:0] s_185;
  wire [16:0] s_186;
  wire [16:0] s_187;
  wire [16:0] s_188;
  wire [12:0] s_189;
  wire [12:0] s_190;
  wire [0:0] s_191;
  wire [12:0] s_192;
  wire [12:0] s_193;
  wire [12:0] s_194;
  wire [12:0] s_195;
  wire [12:0] s_196;
  wire [10:0] s_197;
  wire [10:0] s_198;
  wire [12:0] s_199;
  wire [10:0] s_200;
  wire [10:0] s_201;
  wire [0:0] s_202;
  wire [0:0] s_203;
  wire [12:0] s_204;
  wire [12:0] s_205;
  wire [7:0] s_206;
  wire [7:0] s_207;
  wire [0:0] s_208;
  wire [0:0] s_209;
  wire [6:0] s_210;
  wire [0:0] s_211;
  wire [0:0] s_212;
  wire [5:0] s_213;
  wire [0:0] s_214;
  wire [0:0] s_215;
  wire [4:0] s_216;
  wire [0:0] s_217;
  wire [0:0] s_218;
  wire [3:0] s_219;
  wire [0:0] s_220;
  wire [0:0] s_221;
  wire [2:0] s_222;
  wire [0:0] s_223;
  wire [0:0] s_224;
  wire [1:0] s_225;
  wire [0:0] s_226;
  wire [0:0] s_227;
  wire [0:0] s_228;
  wire [1:0] s_229;
  wire [3:0] s_230;
  wire [7:0] s_231;
  wire [15:0] s_232;
  wire [31:0] s_233;
  wire [63:0] s_234;
  wire [127:0] s_235;
  wire [126:0] s_236;
  wire [125:0] s_237;
  wire [124:0] s_238;
  wire [123:0] s_239;
  wire [122:0] s_240;
  wire [121:0] s_241;
  wire [120:0] s_242;
  wire [119:0] s_243;
  wire [118:0] s_244;
  wire [117:0] s_245;
  wire [116:0] s_246;
  wire [115:0] s_247;
  wire [114:0] s_248;
  wire [113:0] s_249;
  wire [112:0] s_250;
  wire [111:0] s_251;
  wire [110:0] s_252;
  wire [109:0] s_253;
  wire [108:0] s_254;
  wire [107:0] s_255;
  wire [106:0] s_256;
  wire [0:0] s_257;
  wire [0:0] s_258;
  wire [0:0] s_259;
  wire [0:0] s_260;
  wire [0:0] s_261;
  wire [0:0] s_262;
  wire [0:0] s_263;
  wire [0:0] s_264;
  wire [0:0] s_265;
  wire [0:0] s_266;
  wire [0:0] s_267;
  wire [0:0] s_268;
  wire [0:0] s_269;
  wire [0:0] s_270;
  wire [0:0] s_271;
  wire [0:0] s_272;
  wire [0:0] s_273;
  wire [0:0] s_274;
  wire [0:0] s_275;
  wire [0:0] s_276;
  wire [0:0] s_277;
  wire [0:0] s_278;
  wire [0:0] s_279;
  wire [0:0] s_280;
  wire [0:0] s_281;
  wire [0:0] s_282;
  wire [0:0] s_283;
  wire [0:0] s_284;
  wire [0:0] s_285;
  wire [1:0] s_286;
  wire [0:0] s_287;
  wire [0:0] s_288;
  wire [0:0] s_289;
  wire [1:0] s_290;
  wire [0:0] s_291;
  wire [0:0] s_292;
  wire [0:0] s_293;
  wire [0:0] s_294;
  wire [0:0] s_295;
  wire [0:0] s_296;
  wire [1:0] s_297;
  wire [0:0] s_298;
  wire [0:0] s_299;
  wire [0:0] s_300;
  wire [0:0] s_301;
  wire [0:0] s_302;
  wire [0:0] s_303;
  wire [2:0] s_304;
  wire [0:0] s_305;
  wire [0:0] s_306;
  wire [1:0] s_307;
  wire [0:0] s_308;
  wire [0:0] s_309;
  wire [0:0] s_310;
  wire [1:0] s_311;
  wire [3:0] s_312;
  wire [0:0] s_313;
  wire [0:0] s_314;
  wire [0:0] s_315;
  wire [0:0] s_316;
  wire [0:0] s_317;
  wire [0:0] s_318;
  wire [0:0] s_319;
  wire [1:0] s_320;
  wire [0:0] s_321;
  wire [0:0] s_322;
  wire [0:0] s_323;
  wire [1:0] s_324;
  wire [0:0] s_325;
  wire [0:0] s_326;
  wire [0:0] s_327;
  wire [0:0] s_328;
  wire [0:0] s_329;
  wire [0:0] s_330;
  wire [1:0] s_331;
  wire [0:0] s_332;
  wire [0:0] s_333;
  wire [0:0] s_334;
  wire [0:0] s_335;
  wire [0:0] s_336;
  wire [2:0] s_337;
  wire [0:0] s_338;
  wire [0:0] s_339;
  wire [1:0] s_340;
  wire [1:0] s_341;
  wire [1:0] s_342;
  wire [0:0] s_343;
  wire [3:0] s_344;
  wire [0:0] s_345;
  wire [0:0] s_346;
  wire [2:0] s_347;
  wire [0:0] s_348;
  wire [0:0] s_349;
  wire [1:0] s_350;
  wire [0:0] s_351;
  wire [0:0] s_352;
  wire [0:0] s_353;
  wire [1:0] s_354;
  wire [3:0] s_355;
  wire [7:0] s_356;
  wire [0:0] s_357;
  wire [0:0] s_358;
  wire [0:0] s_359;
  wire [0:0] s_360;
  wire [0:0] s_361;
  wire [0:0] s_362;
  wire [0:0] s_363;
  wire [1:0] s_364;
  wire [0:0] s_365;
  wire [0:0] s_366;
  wire [0:0] s_367;
  wire [1:0] s_368;
  wire [0:0] s_369;
  wire [0:0] s_370;
  wire [0:0] s_371;
  wire [0:0] s_372;
  wire [0:0] s_373;
  wire [0:0] s_374;
  wire [1:0] s_375;
  wire [0:0] s_376;
  wire [0:0] s_377;
  wire [0:0] s_378;
  wire [0:0] s_379;
  wire [0:0] s_380;
  wire [0:0] s_381;
  wire [2:0] s_382;
  wire [0:0] s_383;
  wire [0:0] s_384;
  wire [1:0] s_385;
  wire [0:0] s_386;
  wire [0:0] s_387;
  wire [0:0] s_388;
  wire [1:0] s_389;
  wire [3:0] s_390;
  wire [0:0] s_391;
  wire [0:0] s_392;
  wire [0:0] s_393;
  wire [0:0] s_394;
  wire [0:0] s_395;
  wire [0:0] s_396;
  wire [0:0] s_397;
  wire [1:0] s_398;
  wire [0:0] s_399;
  wire [0:0] s_400;
  wire [0:0] s_401;
  wire [1:0] s_402;
  wire [0:0] s_403;
  wire [0:0] s_404;
  wire [0:0] s_405;
  wire [0:0] s_406;
  wire [0:0] s_407;
  wire [0:0] s_408;
  wire [1:0] s_409;
  wire [0:0] s_410;
  wire [0:0] s_411;
  wire [0:0] s_412;
  wire [0:0] s_413;
  wire [0:0] s_414;
  wire [2:0] s_415;
  wire [0:0] s_416;
  wire [0:0] s_417;
  wire [1:0] s_418;
  wire [1:0] s_419;
  wire [1:0] s_420;
  wire [3:0] s_421;
  wire [0:0] s_422;
  wire [0:0] s_423;
  wire [2:0] s_424;
  wire [2:0] s_425;
  wire [2:0] s_426;
  wire [0:0] s_427;
  wire [4:0] s_428;
  wire [0:0] s_429;
  wire [0:0] s_430;
  wire [3:0] s_431;
  wire [0:0] s_432;
  wire [0:0] s_433;
  wire [2:0] s_434;
  wire [0:0] s_435;
  wire [0:0] s_436;
  wire [1:0] s_437;
  wire [0:0] s_438;
  wire [0:0] s_439;
  wire [0:0] s_440;
  wire [1:0] s_441;
  wire [3:0] s_442;
  wire [7:0] s_443;
  wire [15:0] s_444;
  wire [0:0] s_445;
  wire [0:0] s_446;
  wire [0:0] s_447;
  wire [0:0] s_448;
  wire [0:0] s_449;
  wire [0:0] s_450;
  wire [0:0] s_451;
  wire [1:0] s_452;
  wire [0:0] s_453;
  wire [0:0] s_454;
  wire [0:0] s_455;
  wire [1:0] s_456;
  wire [0:0] s_457;
  wire [0:0] s_458;
  wire [0:0] s_459;
  wire [0:0] s_460;
  wire [0:0] s_461;
  wire [0:0] s_462;
  wire [1:0] s_463;
  wire [0:0] s_464;
  wire [0:0] s_465;
  wire [0:0] s_466;
  wire [0:0] s_467;
  wire [0:0] s_468;
  wire [0:0] s_469;
  wire [2:0] s_470;
  wire [0:0] s_471;
  wire [0:0] s_472;
  wire [1:0] s_473;
  wire [0:0] s_474;
  wire [0:0] s_475;
  wire [0:0] s_476;
  wire [1:0] s_477;
  wire [3:0] s_478;
  wire [0:0] s_479;
  wire [0:0] s_480;
  wire [0:0] s_481;
  wire [0:0] s_482;
  wire [0:0] s_483;
  wire [0:0] s_484;
  wire [0:0] s_485;
  wire [1:0] s_486;
  wire [0:0] s_487;
  wire [0:0] s_488;
  wire [0:0] s_489;
  wire [1:0] s_490;
  wire [0:0] s_491;
  wire [0:0] s_492;
  wire [0:0] s_493;
  wire [0:0] s_494;
  wire [0:0] s_495;
  wire [0:0] s_496;
  wire [1:0] s_497;
  wire [0:0] s_498;
  wire [0:0] s_499;
  wire [0:0] s_500;
  wire [0:0] s_501;
  wire [0:0] s_502;
  wire [2:0] s_503;
  wire [0:0] s_504;
  wire [0:0] s_505;
  wire [1:0] s_506;
  wire [1:0] s_507;
  wire [1:0] s_508;
  wire [0:0] s_509;
  wire [3:0] s_510;
  wire [0:0] s_511;
  wire [0:0] s_512;
  wire [2:0] s_513;
  wire [0:0] s_514;
  wire [0:0] s_515;
  wire [1:0] s_516;
  wire [0:0] s_517;
  wire [0:0] s_518;
  wire [0:0] s_519;
  wire [1:0] s_520;
  wire [3:0] s_521;
  wire [7:0] s_522;
  wire [0:0] s_523;
  wire [0:0] s_524;
  wire [0:0] s_525;
  wire [0:0] s_526;
  wire [0:0] s_527;
  wire [0:0] s_528;
  wire [0:0] s_529;
  wire [1:0] s_530;
  wire [0:0] s_531;
  wire [0:0] s_532;
  wire [0:0] s_533;
  wire [1:0] s_534;
  wire [0:0] s_535;
  wire [0:0] s_536;
  wire [0:0] s_537;
  wire [0:0] s_538;
  wire [0:0] s_539;
  wire [0:0] s_540;
  wire [1:0] s_541;
  wire [0:0] s_542;
  wire [0:0] s_543;
  wire [0:0] s_544;
  wire [0:0] s_545;
  wire [0:0] s_546;
  wire [0:0] s_547;
  wire [2:0] s_548;
  wire [0:0] s_549;
  wire [0:0] s_550;
  wire [1:0] s_551;
  wire [0:0] s_552;
  wire [0:0] s_553;
  wire [0:0] s_554;
  wire [1:0] s_555;
  wire [3:0] s_556;
  wire [0:0] s_557;
  wire [0:0] s_558;
  wire [0:0] s_559;
  wire [0:0] s_560;
  wire [0:0] s_561;
  wire [0:0] s_562;
  wire [0:0] s_563;
  wire [1:0] s_564;
  wire [0:0] s_565;
  wire [0:0] s_566;
  wire [0:0] s_567;
  wire [1:0] s_568;
  wire [0:0] s_569;
  wire [0:0] s_570;
  wire [0:0] s_571;
  wire [0:0] s_572;
  wire [0:0] s_573;
  wire [0:0] s_574;
  wire [1:0] s_575;
  wire [0:0] s_576;
  wire [0:0] s_577;
  wire [0:0] s_578;
  wire [0:0] s_579;
  wire [0:0] s_580;
  wire [2:0] s_581;
  wire [0:0] s_582;
  wire [0:0] s_583;
  wire [1:0] s_584;
  wire [1:0] s_585;
  wire [1:0] s_586;
  wire [3:0] s_587;
  wire [0:0] s_588;
  wire [0:0] s_589;
  wire [2:0] s_590;
  wire [2:0] s_591;
  wire [2:0] s_592;
  wire [4:0] s_593;
  wire [0:0] s_594;
  wire [0:0] s_595;
  wire [3:0] s_596;
  wire [3:0] s_597;
  wire [3:0] s_598;
  wire [0:0] s_599;
  wire [5:0] s_600;
  wire [0:0] s_601;
  wire [0:0] s_602;
  wire [4:0] s_603;
  wire [0:0] s_604;
  wire [0:0] s_605;
  wire [3:0] s_606;
  wire [0:0] s_607;
  wire [0:0] s_608;
  wire [2:0] s_609;
  wire [0:0] s_610;
  wire [0:0] s_611;
  wire [1:0] s_612;
  wire [0:0] s_613;
  wire [0:0] s_614;
  wire [0:0] s_615;
  wire [1:0] s_616;
  wire [3:0] s_617;
  wire [7:0] s_618;
  wire [15:0] s_619;
  wire [31:0] s_620;
  wire [0:0] s_621;
  wire [0:0] s_622;
  wire [0:0] s_623;
  wire [0:0] s_624;
  wire [0:0] s_625;
  wire [0:0] s_626;
  wire [0:0] s_627;
  wire [1:0] s_628;
  wire [0:0] s_629;
  wire [0:0] s_630;
  wire [0:0] s_631;
  wire [1:0] s_632;
  wire [0:0] s_633;
  wire [0:0] s_634;
  wire [0:0] s_635;
  wire [0:0] s_636;
  wire [0:0] s_637;
  wire [0:0] s_638;
  wire [1:0] s_639;
  wire [0:0] s_640;
  wire [0:0] s_641;
  wire [0:0] s_642;
  wire [0:0] s_643;
  wire [0:0] s_644;
  wire [0:0] s_645;
  wire [2:0] s_646;
  wire [0:0] s_647;
  wire [0:0] s_648;
  wire [1:0] s_649;
  wire [0:0] s_650;
  wire [0:0] s_651;
  wire [0:0] s_652;
  wire [1:0] s_653;
  wire [3:0] s_654;
  wire [0:0] s_655;
  wire [0:0] s_656;
  wire [0:0] s_657;
  wire [0:0] s_658;
  wire [0:0] s_659;
  wire [0:0] s_660;
  wire [0:0] s_661;
  wire [1:0] s_662;
  wire [0:0] s_663;
  wire [0:0] s_664;
  wire [0:0] s_665;
  wire [1:0] s_666;
  wire [0:0] s_667;
  wire [0:0] s_668;
  wire [0:0] s_669;
  wire [0:0] s_670;
  wire [0:0] s_671;
  wire [0:0] s_672;
  wire [1:0] s_673;
  wire [0:0] s_674;
  wire [0:0] s_675;
  wire [0:0] s_676;
  wire [0:0] s_677;
  wire [0:0] s_678;
  wire [2:0] s_679;
  wire [0:0] s_680;
  wire [0:0] s_681;
  wire [1:0] s_682;
  wire [1:0] s_683;
  wire [1:0] s_684;
  wire [0:0] s_685;
  wire [3:0] s_686;
  wire [0:0] s_687;
  wire [0:0] s_688;
  wire [2:0] s_689;
  wire [0:0] s_690;
  wire [0:0] s_691;
  wire [1:0] s_692;
  wire [0:0] s_693;
  wire [0:0] s_694;
  wire [0:0] s_695;
  wire [1:0] s_696;
  wire [3:0] s_697;
  wire [7:0] s_698;
  wire [0:0] s_699;
  wire [0:0] s_700;
  wire [0:0] s_701;
  wire [0:0] s_702;
  wire [0:0] s_703;
  wire [0:0] s_704;
  wire [0:0] s_705;
  wire [1:0] s_706;
  wire [0:0] s_707;
  wire [0:0] s_708;
  wire [0:0] s_709;
  wire [1:0] s_710;
  wire [0:0] s_711;
  wire [0:0] s_712;
  wire [0:0] s_713;
  wire [0:0] s_714;
  wire [0:0] s_715;
  wire [0:0] s_716;
  wire [1:0] s_717;
  wire [0:0] s_718;
  wire [0:0] s_719;
  wire [0:0] s_720;
  wire [0:0] s_721;
  wire [0:0] s_722;
  wire [0:0] s_723;
  wire [2:0] s_724;
  wire [0:0] s_725;
  wire [0:0] s_726;
  wire [1:0] s_727;
  wire [0:0] s_728;
  wire [0:0] s_729;
  wire [0:0] s_730;
  wire [1:0] s_731;
  wire [3:0] s_732;
  wire [0:0] s_733;
  wire [0:0] s_734;
  wire [0:0] s_735;
  wire [0:0] s_736;
  wire [0:0] s_737;
  wire [0:0] s_738;
  wire [0:0] s_739;
  wire [1:0] s_740;
  wire [0:0] s_741;
  wire [0:0] s_742;
  wire [0:0] s_743;
  wire [1:0] s_744;
  wire [0:0] s_745;
  wire [0:0] s_746;
  wire [0:0] s_747;
  wire [0:0] s_748;
  wire [0:0] s_749;
  wire [0:0] s_750;
  wire [1:0] s_751;
  wire [0:0] s_752;
  wire [0:0] s_753;
  wire [0:0] s_754;
  wire [0:0] s_755;
  wire [0:0] s_756;
  wire [2:0] s_757;
  wire [0:0] s_758;
  wire [0:0] s_759;
  wire [1:0] s_760;
  wire [1:0] s_761;
  wire [1:0] s_762;
  wire [3:0] s_763;
  wire [0:0] s_764;
  wire [0:0] s_765;
  wire [2:0] s_766;
  wire [2:0] s_767;
  wire [2:0] s_768;
  wire [0:0] s_769;
  wire [4:0] s_770;
  wire [0:0] s_771;
  wire [0:0] s_772;
  wire [3:0] s_773;
  wire [0:0] s_774;
  wire [0:0] s_775;
  wire [2:0] s_776;
  wire [0:0] s_777;
  wire [0:0] s_778;
  wire [1:0] s_779;
  wire [0:0] s_780;
  wire [0:0] s_781;
  wire [0:0] s_782;
  wire [1:0] s_783;
  wire [3:0] s_784;
  wire [7:0] s_785;
  wire [15:0] s_786;
  wire [0:0] s_787;
  wire [0:0] s_788;
  wire [0:0] s_789;
  wire [0:0] s_790;
  wire [0:0] s_791;
  wire [0:0] s_792;
  wire [0:0] s_793;
  wire [1:0] s_794;
  wire [0:0] s_795;
  wire [0:0] s_796;
  wire [0:0] s_797;
  wire [1:0] s_798;
  wire [0:0] s_799;
  wire [0:0] s_800;
  wire [0:0] s_801;
  wire [0:0] s_802;
  wire [0:0] s_803;
  wire [0:0] s_804;
  wire [1:0] s_805;
  wire [0:0] s_806;
  wire [0:0] s_807;
  wire [0:0] s_808;
  wire [0:0] s_809;
  wire [0:0] s_810;
  wire [0:0] s_811;
  wire [2:0] s_812;
  wire [0:0] s_813;
  wire [0:0] s_814;
  wire [1:0] s_815;
  wire [0:0] s_816;
  wire [0:0] s_817;
  wire [0:0] s_818;
  wire [1:0] s_819;
  wire [3:0] s_820;
  wire [0:0] s_821;
  wire [0:0] s_822;
  wire [0:0] s_823;
  wire [0:0] s_824;
  wire [0:0] s_825;
  wire [0:0] s_826;
  wire [0:0] s_827;
  wire [1:0] s_828;
  wire [0:0] s_829;
  wire [0:0] s_830;
  wire [0:0] s_831;
  wire [1:0] s_832;
  wire [0:0] s_833;
  wire [0:0] s_834;
  wire [0:0] s_835;
  wire [0:0] s_836;
  wire [0:0] s_837;
  wire [0:0] s_838;
  wire [1:0] s_839;
  wire [0:0] s_840;
  wire [0:0] s_841;
  wire [0:0] s_842;
  wire [0:0] s_843;
  wire [0:0] s_844;
  wire [2:0] s_845;
  wire [0:0] s_846;
  wire [0:0] s_847;
  wire [1:0] s_848;
  wire [1:0] s_849;
  wire [1:0] s_850;
  wire [0:0] s_851;
  wire [3:0] s_852;
  wire [0:0] s_853;
  wire [0:0] s_854;
  wire [2:0] s_855;
  wire [0:0] s_856;
  wire [0:0] s_857;
  wire [1:0] s_858;
  wire [0:0] s_859;
  wire [0:0] s_860;
  wire [0:0] s_861;
  wire [1:0] s_862;
  wire [3:0] s_863;
  wire [7:0] s_864;
  wire [0:0] s_865;
  wire [0:0] s_866;
  wire [0:0] s_867;
  wire [0:0] s_868;
  wire [0:0] s_869;
  wire [0:0] s_870;
  wire [0:0] s_871;
  wire [1:0] s_872;
  wire [0:0] s_873;
  wire [0:0] s_874;
  wire [0:0] s_875;
  wire [1:0] s_876;
  wire [0:0] s_877;
  wire [0:0] s_878;
  wire [0:0] s_879;
  wire [0:0] s_880;
  wire [0:0] s_881;
  wire [0:0] s_882;
  wire [1:0] s_883;
  wire [0:0] s_884;
  wire [0:0] s_885;
  wire [0:0] s_886;
  wire [0:0] s_887;
  wire [0:0] s_888;
  wire [0:0] s_889;
  wire [2:0] s_890;
  wire [0:0] s_891;
  wire [0:0] s_892;
  wire [1:0] s_893;
  wire [0:0] s_894;
  wire [0:0] s_895;
  wire [0:0] s_896;
  wire [1:0] s_897;
  wire [3:0] s_898;
  wire [0:0] s_899;
  wire [0:0] s_900;
  wire [0:0] s_901;
  wire [0:0] s_902;
  wire [0:0] s_903;
  wire [0:0] s_904;
  wire [0:0] s_905;
  wire [1:0] s_906;
  wire [0:0] s_907;
  wire [0:0] s_908;
  wire [0:0] s_909;
  wire [1:0] s_910;
  wire [0:0] s_911;
  wire [0:0] s_912;
  wire [0:0] s_913;
  wire [0:0] s_914;
  wire [0:0] s_915;
  wire [0:0] s_916;
  wire [1:0] s_917;
  wire [0:0] s_918;
  wire [0:0] s_919;
  wire [0:0] s_920;
  wire [0:0] s_921;
  wire [0:0] s_922;
  wire [2:0] s_923;
  wire [0:0] s_924;
  wire [0:0] s_925;
  wire [1:0] s_926;
  wire [1:0] s_927;
  wire [1:0] s_928;
  wire [3:0] s_929;
  wire [0:0] s_930;
  wire [0:0] s_931;
  wire [2:0] s_932;
  wire [2:0] s_933;
  wire [2:0] s_934;
  wire [4:0] s_935;
  wire [0:0] s_936;
  wire [0:0] s_937;
  wire [3:0] s_938;
  wire [3:0] s_939;
  wire [3:0] s_940;
  wire [5:0] s_941;
  wire [0:0] s_942;
  wire [0:0] s_943;
  wire [4:0] s_944;
  wire [4:0] s_945;
  wire [4:0] s_946;
  wire [0:0] s_947;
  wire [6:0] s_948;
  wire [0:0] s_949;
  wire [0:0] s_950;
  wire [5:0] s_951;
  wire [0:0] s_952;
  wire [0:0] s_953;
  wire [4:0] s_954;
  wire [0:0] s_955;
  wire [0:0] s_956;
  wire [3:0] s_957;
  wire [0:0] s_958;
  wire [0:0] s_959;
  wire [2:0] s_960;
  wire [0:0] s_961;
  wire [0:0] s_962;
  wire [1:0] s_963;
  wire [0:0] s_964;
  wire [0:0] s_965;
  wire [0:0] s_966;
  wire [1:0] s_967;
  wire [3:0] s_968;
  wire [7:0] s_969;
  wire [15:0] s_970;
  wire [31:0] s_971;
  wire [63:0] s_972;
  wire [0:0] s_973;
  wire [0:0] s_974;
  wire [0:0] s_975;
  wire [0:0] s_976;
  wire [0:0] s_977;
  wire [0:0] s_978;
  wire [0:0] s_979;
  wire [1:0] s_980;
  wire [0:0] s_981;
  wire [0:0] s_982;
  wire [0:0] s_983;
  wire [1:0] s_984;
  wire [0:0] s_985;
  wire [0:0] s_986;
  wire [0:0] s_987;
  wire [0:0] s_988;
  wire [0:0] s_989;
  wire [0:0] s_990;
  wire [1:0] s_991;
  wire [0:0] s_992;
  wire [0:0] s_993;
  wire [0:0] s_994;
  wire [0:0] s_995;
  wire [0:0] s_996;
  wire [0:0] s_997;
  wire [2:0] s_998;
  wire [0:0] s_999;
  wire [0:0] s_1000;
  wire [1:0] s_1001;
  wire [0:0] s_1002;
  wire [0:0] s_1003;
  wire [0:0] s_1004;
  wire [1:0] s_1005;
  wire [3:0] s_1006;
  wire [0:0] s_1007;
  wire [0:0] s_1008;
  wire [0:0] s_1009;
  wire [0:0] s_1010;
  wire [0:0] s_1011;
  wire [0:0] s_1012;
  wire [0:0] s_1013;
  wire [1:0] s_1014;
  wire [0:0] s_1015;
  wire [0:0] s_1016;
  wire [0:0] s_1017;
  wire [1:0] s_1018;
  wire [0:0] s_1019;
  wire [0:0] s_1020;
  wire [0:0] s_1021;
  wire [0:0] s_1022;
  wire [0:0] s_1023;
  wire [0:0] s_1024;
  wire [1:0] s_1025;
  wire [0:0] s_1026;
  wire [0:0] s_1027;
  wire [0:0] s_1028;
  wire [0:0] s_1029;
  wire [0:0] s_1030;
  wire [2:0] s_1031;
  wire [0:0] s_1032;
  wire [0:0] s_1033;
  wire [1:0] s_1034;
  wire [1:0] s_1035;
  wire [1:0] s_1036;
  wire [0:0] s_1037;
  wire [3:0] s_1038;
  wire [0:0] s_1039;
  wire [0:0] s_1040;
  wire [2:0] s_1041;
  wire [0:0] s_1042;
  wire [0:0] s_1043;
  wire [1:0] s_1044;
  wire [0:0] s_1045;
  wire [0:0] s_1046;
  wire [0:0] s_1047;
  wire [1:0] s_1048;
  wire [3:0] s_1049;
  wire [7:0] s_1050;
  wire [0:0] s_1051;
  wire [0:0] s_1052;
  wire [0:0] s_1053;
  wire [0:0] s_1054;
  wire [0:0] s_1055;
  wire [0:0] s_1056;
  wire [0:0] s_1057;
  wire [1:0] s_1058;
  wire [0:0] s_1059;
  wire [0:0] s_1060;
  wire [0:0] s_1061;
  wire [1:0] s_1062;
  wire [0:0] s_1063;
  wire [0:0] s_1064;
  wire [0:0] s_1065;
  wire [0:0] s_1066;
  wire [0:0] s_1067;
  wire [0:0] s_1068;
  wire [1:0] s_1069;
  wire [0:0] s_1070;
  wire [0:0] s_1071;
  wire [0:0] s_1072;
  wire [0:0] s_1073;
  wire [0:0] s_1074;
  wire [0:0] s_1075;
  wire [2:0] s_1076;
  wire [0:0] s_1077;
  wire [0:0] s_1078;
  wire [1:0] s_1079;
  wire [0:0] s_1080;
  wire [0:0] s_1081;
  wire [0:0] s_1082;
  wire [1:0] s_1083;
  wire [3:0] s_1084;
  wire [0:0] s_1085;
  wire [0:0] s_1086;
  wire [0:0] s_1087;
  wire [0:0] s_1088;
  wire [0:0] s_1089;
  wire [0:0] s_1090;
  wire [0:0] s_1091;
  wire [1:0] s_1092;
  wire [0:0] s_1093;
  wire [0:0] s_1094;
  wire [0:0] s_1095;
  wire [1:0] s_1096;
  wire [0:0] s_1097;
  wire [0:0] s_1098;
  wire [0:0] s_1099;
  wire [0:0] s_1100;
  wire [0:0] s_1101;
  wire [0:0] s_1102;
  wire [1:0] s_1103;
  wire [0:0] s_1104;
  wire [0:0] s_1105;
  wire [0:0] s_1106;
  wire [0:0] s_1107;
  wire [0:0] s_1108;
  wire [2:0] s_1109;
  wire [0:0] s_1110;
  wire [0:0] s_1111;
  wire [1:0] s_1112;
  wire [1:0] s_1113;
  wire [1:0] s_1114;
  wire [3:0] s_1115;
  wire [0:0] s_1116;
  wire [0:0] s_1117;
  wire [2:0] s_1118;
  wire [2:0] s_1119;
  wire [2:0] s_1120;
  wire [0:0] s_1121;
  wire [4:0] s_1122;
  wire [0:0] s_1123;
  wire [0:0] s_1124;
  wire [3:0] s_1125;
  wire [0:0] s_1126;
  wire [0:0] s_1127;
  wire [2:0] s_1128;
  wire [0:0] s_1129;
  wire [0:0] s_1130;
  wire [1:0] s_1131;
  wire [0:0] s_1132;
  wire [0:0] s_1133;
  wire [0:0] s_1134;
  wire [1:0] s_1135;
  wire [3:0] s_1136;
  wire [7:0] s_1137;
  wire [15:0] s_1138;
  wire [0:0] s_1139;
  wire [0:0] s_1140;
  wire [0:0] s_1141;
  wire [0:0] s_1142;
  wire [0:0] s_1143;
  wire [0:0] s_1144;
  wire [0:0] s_1145;
  wire [1:0] s_1146;
  wire [0:0] s_1147;
  wire [0:0] s_1148;
  wire [0:0] s_1149;
  wire [1:0] s_1150;
  wire [0:0] s_1151;
  wire [0:0] s_1152;
  wire [0:0] s_1153;
  wire [0:0] s_1154;
  wire [0:0] s_1155;
  wire [0:0] s_1156;
  wire [1:0] s_1157;
  wire [0:0] s_1158;
  wire [0:0] s_1159;
  wire [0:0] s_1160;
  wire [0:0] s_1161;
  wire [0:0] s_1162;
  wire [0:0] s_1163;
  wire [2:0] s_1164;
  wire [0:0] s_1165;
  wire [0:0] s_1166;
  wire [1:0] s_1167;
  wire [0:0] s_1168;
  wire [0:0] s_1169;
  wire [0:0] s_1170;
  wire [1:0] s_1171;
  wire [3:0] s_1172;
  wire [0:0] s_1173;
  wire [0:0] s_1174;
  wire [0:0] s_1175;
  wire [0:0] s_1176;
  wire [0:0] s_1177;
  wire [0:0] s_1178;
  wire [0:0] s_1179;
  wire [1:0] s_1180;
  wire [0:0] s_1181;
  wire [0:0] s_1182;
  wire [0:0] s_1183;
  wire [1:0] s_1184;
  wire [0:0] s_1185;
  wire [0:0] s_1186;
  wire [0:0] s_1187;
  wire [0:0] s_1188;
  wire [0:0] s_1189;
  wire [0:0] s_1190;
  wire [1:0] s_1191;
  wire [0:0] s_1192;
  wire [0:0] s_1193;
  wire [0:0] s_1194;
  wire [0:0] s_1195;
  wire [0:0] s_1196;
  wire [2:0] s_1197;
  wire [0:0] s_1198;
  wire [0:0] s_1199;
  wire [1:0] s_1200;
  wire [1:0] s_1201;
  wire [1:0] s_1202;
  wire [0:0] s_1203;
  wire [3:0] s_1204;
  wire [0:0] s_1205;
  wire [0:0] s_1206;
  wire [2:0] s_1207;
  wire [0:0] s_1208;
  wire [0:0] s_1209;
  wire [1:0] s_1210;
  wire [0:0] s_1211;
  wire [0:0] s_1212;
  wire [0:0] s_1213;
  wire [1:0] s_1214;
  wire [3:0] s_1215;
  wire [7:0] s_1216;
  wire [0:0] s_1217;
  wire [0:0] s_1218;
  wire [0:0] s_1219;
  wire [0:0] s_1220;
  wire [0:0] s_1221;
  wire [0:0] s_1222;
  wire [0:0] s_1223;
  wire [1:0] s_1224;
  wire [0:0] s_1225;
  wire [0:0] s_1226;
  wire [0:0] s_1227;
  wire [1:0] s_1228;
  wire [0:0] s_1229;
  wire [0:0] s_1230;
  wire [0:0] s_1231;
  wire [0:0] s_1232;
  wire [0:0] s_1233;
  wire [0:0] s_1234;
  wire [1:0] s_1235;
  wire [0:0] s_1236;
  wire [0:0] s_1237;
  wire [0:0] s_1238;
  wire [0:0] s_1239;
  wire [0:0] s_1240;
  wire [0:0] s_1241;
  wire [2:0] s_1242;
  wire [0:0] s_1243;
  wire [0:0] s_1244;
  wire [1:0] s_1245;
  wire [0:0] s_1246;
  wire [0:0] s_1247;
  wire [0:0] s_1248;
  wire [1:0] s_1249;
  wire [3:0] s_1250;
  wire [0:0] s_1251;
  wire [0:0] s_1252;
  wire [0:0] s_1253;
  wire [0:0] s_1254;
  wire [0:0] s_1255;
  wire [0:0] s_1256;
  wire [0:0] s_1257;
  wire [1:0] s_1258;
  wire [0:0] s_1259;
  wire [0:0] s_1260;
  wire [0:0] s_1261;
  wire [1:0] s_1262;
  wire [0:0] s_1263;
  wire [0:0] s_1264;
  wire [0:0] s_1265;
  wire [0:0] s_1266;
  wire [0:0] s_1267;
  wire [0:0] s_1268;
  wire [1:0] s_1269;
  wire [0:0] s_1270;
  wire [0:0] s_1271;
  wire [0:0] s_1272;
  wire [0:0] s_1273;
  wire [0:0] s_1274;
  wire [2:0] s_1275;
  wire [0:0] s_1276;
  wire [0:0] s_1277;
  wire [1:0] s_1278;
  wire [1:0] s_1279;
  wire [1:0] s_1280;
  wire [3:0] s_1281;
  wire [0:0] s_1282;
  wire [0:0] s_1283;
  wire [2:0] s_1284;
  wire [2:0] s_1285;
  wire [2:0] s_1286;
  wire [4:0] s_1287;
  wire [0:0] s_1288;
  wire [0:0] s_1289;
  wire [3:0] s_1290;
  wire [3:0] s_1291;
  wire [3:0] s_1292;
  wire [0:0] s_1293;
  wire [5:0] s_1294;
  wire [0:0] s_1295;
  wire [0:0] s_1296;
  wire [4:0] s_1297;
  wire [0:0] s_1298;
  wire [0:0] s_1299;
  wire [3:0] s_1300;
  wire [0:0] s_1301;
  wire [0:0] s_1302;
  wire [2:0] s_1303;
  wire [0:0] s_1304;
  wire [0:0] s_1305;
  wire [1:0] s_1306;
  wire [0:0] s_1307;
  wire [0:0] s_1308;
  wire [0:0] s_1309;
  wire [1:0] s_1310;
  wire [3:0] s_1311;
  wire [7:0] s_1312;
  wire [15:0] s_1313;
  wire [31:0] s_1314;
  wire [0:0] s_1315;
  wire [0:0] s_1316;
  wire [0:0] s_1317;
  wire [0:0] s_1318;
  wire [0:0] s_1319;
  wire [0:0] s_1320;
  wire [0:0] s_1321;
  wire [1:0] s_1322;
  wire [0:0] s_1323;
  wire [0:0] s_1324;
  wire [0:0] s_1325;
  wire [1:0] s_1326;
  wire [0:0] s_1327;
  wire [0:0] s_1328;
  wire [0:0] s_1329;
  wire [0:0] s_1330;
  wire [0:0] s_1331;
  wire [0:0] s_1332;
  wire [1:0] s_1333;
  wire [0:0] s_1334;
  wire [0:0] s_1335;
  wire [0:0] s_1336;
  wire [0:0] s_1337;
  wire [0:0] s_1338;
  wire [0:0] s_1339;
  wire [2:0] s_1340;
  wire [0:0] s_1341;
  wire [0:0] s_1342;
  wire [1:0] s_1343;
  wire [0:0] s_1344;
  wire [0:0] s_1345;
  wire [0:0] s_1346;
  wire [1:0] s_1347;
  wire [3:0] s_1348;
  wire [0:0] s_1349;
  wire [0:0] s_1350;
  wire [0:0] s_1351;
  wire [0:0] s_1352;
  wire [0:0] s_1353;
  wire [0:0] s_1354;
  wire [0:0] s_1355;
  wire [1:0] s_1356;
  wire [0:0] s_1357;
  wire [0:0] s_1358;
  wire [0:0] s_1359;
  wire [1:0] s_1360;
  wire [0:0] s_1361;
  wire [0:0] s_1362;
  wire [0:0] s_1363;
  wire [0:0] s_1364;
  wire [0:0] s_1365;
  wire [0:0] s_1366;
  wire [1:0] s_1367;
  wire [0:0] s_1368;
  wire [0:0] s_1369;
  wire [0:0] s_1370;
  wire [0:0] s_1371;
  wire [0:0] s_1372;
  wire [2:0] s_1373;
  wire [0:0] s_1374;
  wire [0:0] s_1375;
  wire [1:0] s_1376;
  wire [1:0] s_1377;
  wire [1:0] s_1378;
  wire [0:0] s_1379;
  wire [3:0] s_1380;
  wire [0:0] s_1381;
  wire [0:0] s_1382;
  wire [2:0] s_1383;
  wire [0:0] s_1384;
  wire [0:0] s_1385;
  wire [1:0] s_1386;
  wire [0:0] s_1387;
  wire [0:0] s_1388;
  wire [0:0] s_1389;
  wire [1:0] s_1390;
  wire [3:0] s_1391;
  wire [7:0] s_1392;
  wire [0:0] s_1393;
  wire [0:0] s_1394;
  wire [0:0] s_1395;
  wire [0:0] s_1396;
  wire [0:0] s_1397;
  wire [0:0] s_1398;
  wire [0:0] s_1399;
  wire [1:0] s_1400;
  wire [0:0] s_1401;
  wire [0:0] s_1402;
  wire [0:0] s_1403;
  wire [1:0] s_1404;
  wire [0:0] s_1405;
  wire [0:0] s_1406;
  wire [0:0] s_1407;
  wire [0:0] s_1408;
  wire [0:0] s_1409;
  wire [0:0] s_1410;
  wire [1:0] s_1411;
  wire [0:0] s_1412;
  wire [0:0] s_1413;
  wire [0:0] s_1414;
  wire [0:0] s_1415;
  wire [0:0] s_1416;
  wire [0:0] s_1417;
  wire [2:0] s_1418;
  wire [0:0] s_1419;
  wire [0:0] s_1420;
  wire [1:0] s_1421;
  wire [0:0] s_1422;
  wire [0:0] s_1423;
  wire [0:0] s_1424;
  wire [1:0] s_1425;
  wire [3:0] s_1426;
  wire [0:0] s_1427;
  wire [0:0] s_1428;
  wire [0:0] s_1429;
  wire [0:0] s_1430;
  wire [0:0] s_1431;
  wire [0:0] s_1432;
  wire [0:0] s_1433;
  wire [1:0] s_1434;
  wire [0:0] s_1435;
  wire [0:0] s_1436;
  wire [0:0] s_1437;
  wire [1:0] s_1438;
  wire [0:0] s_1439;
  wire [0:0] s_1440;
  wire [0:0] s_1441;
  wire [0:0] s_1442;
  wire [0:0] s_1443;
  wire [0:0] s_1444;
  wire [1:0] s_1445;
  wire [0:0] s_1446;
  wire [0:0] s_1447;
  wire [0:0] s_1448;
  wire [0:0] s_1449;
  wire [0:0] s_1450;
  wire [2:0] s_1451;
  wire [0:0] s_1452;
  wire [0:0] s_1453;
  wire [1:0] s_1454;
  wire [1:0] s_1455;
  wire [1:0] s_1456;
  wire [3:0] s_1457;
  wire [0:0] s_1458;
  wire [0:0] s_1459;
  wire [2:0] s_1460;
  wire [2:0] s_1461;
  wire [2:0] s_1462;
  wire [0:0] s_1463;
  wire [4:0] s_1464;
  wire [0:0] s_1465;
  wire [0:0] s_1466;
  wire [3:0] s_1467;
  wire [0:0] s_1468;
  wire [0:0] s_1469;
  wire [2:0] s_1470;
  wire [0:0] s_1471;
  wire [0:0] s_1472;
  wire [1:0] s_1473;
  wire [0:0] s_1474;
  wire [0:0] s_1475;
  wire [0:0] s_1476;
  wire [1:0] s_1477;
  wire [3:0] s_1478;
  wire [7:0] s_1479;
  wire [15:0] s_1480;
  wire [0:0] s_1481;
  wire [0:0] s_1482;
  wire [0:0] s_1483;
  wire [0:0] s_1484;
  wire [0:0] s_1485;
  wire [0:0] s_1486;
  wire [0:0] s_1487;
  wire [1:0] s_1488;
  wire [0:0] s_1489;
  wire [0:0] s_1490;
  wire [0:0] s_1491;
  wire [1:0] s_1492;
  wire [0:0] s_1493;
  wire [0:0] s_1494;
  wire [0:0] s_1495;
  wire [0:0] s_1496;
  wire [0:0] s_1497;
  wire [0:0] s_1498;
  wire [1:0] s_1499;
  wire [0:0] s_1500;
  wire [0:0] s_1501;
  wire [0:0] s_1502;
  wire [0:0] s_1503;
  wire [0:0] s_1504;
  wire [0:0] s_1505;
  wire [2:0] s_1506;
  wire [0:0] s_1507;
  wire [0:0] s_1508;
  wire [1:0] s_1509;
  wire [0:0] s_1510;
  wire [0:0] s_1511;
  wire [0:0] s_1512;
  wire [1:0] s_1513;
  wire [3:0] s_1514;
  wire [0:0] s_1515;
  wire [0:0] s_1516;
  wire [0:0] s_1517;
  wire [0:0] s_1518;
  wire [0:0] s_1519;
  wire [0:0] s_1520;
  wire [0:0] s_1521;
  wire [1:0] s_1522;
  wire [0:0] s_1523;
  wire [0:0] s_1524;
  wire [0:0] s_1525;
  wire [1:0] s_1526;
  wire [0:0] s_1527;
  wire [0:0] s_1528;
  wire [0:0] s_1529;
  wire [0:0] s_1530;
  wire [0:0] s_1531;
  wire [0:0] s_1532;
  wire [1:0] s_1533;
  wire [0:0] s_1534;
  wire [0:0] s_1535;
  wire [0:0] s_1536;
  wire [0:0] s_1537;
  wire [0:0] s_1538;
  wire [2:0] s_1539;
  wire [0:0] s_1540;
  wire [0:0] s_1541;
  wire [1:0] s_1542;
  wire [1:0] s_1543;
  wire [1:0] s_1544;
  wire [0:0] s_1545;
  wire [3:0] s_1546;
  wire [0:0] s_1547;
  wire [0:0] s_1548;
  wire [2:0] s_1549;
  wire [0:0] s_1550;
  wire [0:0] s_1551;
  wire [1:0] s_1552;
  wire [0:0] s_1553;
  wire [0:0] s_1554;
  wire [0:0] s_1555;
  wire [1:0] s_1556;
  wire [3:0] s_1557;
  wire [7:0] s_1558;
  wire [0:0] s_1559;
  wire [0:0] s_1560;
  wire [0:0] s_1561;
  wire [0:0] s_1562;
  wire [0:0] s_1563;
  wire [0:0] s_1564;
  wire [0:0] s_1565;
  wire [1:0] s_1566;
  wire [0:0] s_1567;
  wire [0:0] s_1568;
  wire [0:0] s_1569;
  wire [1:0] s_1570;
  wire [0:0] s_1571;
  wire [0:0] s_1572;
  wire [0:0] s_1573;
  wire [0:0] s_1574;
  wire [0:0] s_1575;
  wire [0:0] s_1576;
  wire [1:0] s_1577;
  wire [0:0] s_1578;
  wire [0:0] s_1579;
  wire [0:0] s_1580;
  wire [0:0] s_1581;
  wire [0:0] s_1582;
  wire [0:0] s_1583;
  wire [2:0] s_1584;
  wire [0:0] s_1585;
  wire [0:0] s_1586;
  wire [1:0] s_1587;
  wire [0:0] s_1588;
  wire [0:0] s_1589;
  wire [0:0] s_1590;
  wire [1:0] s_1591;
  wire [3:0] s_1592;
  wire [0:0] s_1593;
  wire [0:0] s_1594;
  wire [0:0] s_1595;
  wire [0:0] s_1596;
  wire [0:0] s_1597;
  wire [0:0] s_1598;
  wire [0:0] s_1599;
  wire [1:0] s_1600;
  wire [0:0] s_1601;
  wire [0:0] s_1602;
  wire [0:0] s_1603;
  wire [1:0] s_1604;
  wire [0:0] s_1605;
  wire [0:0] s_1606;
  wire [0:0] s_1607;
  wire [0:0] s_1608;
  wire [0:0] s_1609;
  wire [0:0] s_1610;
  wire [1:0] s_1611;
  wire [0:0] s_1612;
  wire [0:0] s_1613;
  wire [0:0] s_1614;
  wire [0:0] s_1615;
  wire [0:0] s_1616;
  wire [2:0] s_1617;
  wire [0:0] s_1618;
  wire [0:0] s_1619;
  wire [1:0] s_1620;
  wire [1:0] s_1621;
  wire [1:0] s_1622;
  wire [3:0] s_1623;
  wire [0:0] s_1624;
  wire [0:0] s_1625;
  wire [2:0] s_1626;
  wire [2:0] s_1627;
  wire [2:0] s_1628;
  wire [4:0] s_1629;
  wire [0:0] s_1630;
  wire [0:0] s_1631;
  wire [3:0] s_1632;
  wire [3:0] s_1633;
  wire [3:0] s_1634;
  wire [5:0] s_1635;
  wire [0:0] s_1636;
  wire [0:0] s_1637;
  wire [4:0] s_1638;
  wire [4:0] s_1639;
  wire [4:0] s_1640;
  wire [6:0] s_1641;
  wire [0:0] s_1642;
  wire [0:0] s_1643;
  wire [5:0] s_1644;
  wire [5:0] s_1645;
  wire [5:0] s_1646;
  wire [12:0] s_1647;
  wire [12:0] s_1648;
  wire [12:0] s_1649;
  wire [12:0] s_1650;
  wire [12:0] s_1651;
  wire [0:0] s_1652;
  wire [12:0] s_1653;
  wire [12:0] s_1654;
  wire [0:0] s_1655;
  wire [52:0] s_1656;
  wire [0:0] s_1657;
  wire [0:0] s_1658;
  wire [0:0] s_1659;
  wire [0:0] s_1660;
  wire [0:0] s_1661;
  wire [0:0] s_1662;
  wire [0:0] s_1663;
  wire [0:0] s_1664;
  wire [0:0] s_1665;
  wire [50:0] s_1666;
  wire [52:0] s_1667;
  wire [0:0] s_1668;
  wire [0:0] s_1669;
  wire [52:0] s_1670;
  wire [0:0] s_1671;
  wire [63:0] s_1672;
  wire [11:0] s_1673;
  wire [0:0] s_1674;
  wire [10:0] s_1675;
  wire [10:0] s_1676;
  wire [12:0] s_1677;
  wire [12:0] s_1678;
  wire [12:0] s_1679;
  wire [12:0] s_1680;
  wire [12:0] s_1681;
  wire [12:0] s_1682;
  wire [9:0] s_1683;
  wire [51:0] s_1684;
  wire [0:0] s_1685;
  wire [0:0] s_1686;
  wire [10:0] s_1687;
  wire [0:0] s_1688;
  wire [0:0] s_1689;
  wire [0:0] s_1690;
  wire [52:0] s_1691;
  wire [0:0] s_1692;
  wire [0:0] s_1693;
  wire [0:0] s_1694;
  wire [11:0] s_1695;
  wire [0:0] s_1696;
  wire [0:0] s_1697;
  wire [0:0] s_1698;
  wire [10:0] s_1699;
  wire [0:0] s_1700;
  wire [51:0] s_1701;
  wire [0:0] s_1702;
  wire [0:0] s_1703;
  wire [0:0] s_1704;
  wire [10:0] s_1705;
  wire [0:0] s_1706;
  wire [51:0] s_1707;
  wire [0:0] s_1708;
  wire [0:0] s_1709;
  wire [0:0] s_1710;
  wire [0:0] s_1711;
  wire [10:0] s_1712;
  wire [0:0] s_1713;
  wire [51:0] s_1714;
  wire [0:0] s_1715;
  wire [0:0] s_1716;
  wire [10:0] s_1717;
  wire [0:0] s_1718;
  wire [51:0] s_1719;

  assign s_0 = s_1708?s_1:s_9;
  dq #(64, 21) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_8};
  assign s_3 = s_4 ^ s_6;
  assign s_4 = s_5[63];
  assign s_5 = double_mul_a;
  assign s_6 = s_7[63];
  assign s_7 = double_mul_b;
  assign s_8 = 63'd9221120237041090560;
  assign s_9 = s_1692?s_10:s_13;
  dq #(64, 21) dq_s_10 (clk, s_10, s_11);
  assign s_11 = {s_3,s_12};
  assign s_12 = 63'd9218868437227405312;
  assign s_13 = s_1690?s_14:s_17;
  dq #(64, 21) dq_s_14 (clk, s_14, s_15);
  assign s_15 = {s_3,s_16};
  assign s_16 = 63'd0;
  assign s_17 = s_1685?s_18:s_1672;
  assign s_18 = {s_19,s_22};
  dq #(12, 21) dq_s_19 (clk, s_19, s_20);
  assign s_20 = {s_3,s_21};
  assign s_21 = 11'd0;
  assign s_22 = s_23[51:0];
  dq #(53, 1) dq_s_23 (clk, s_23, s_24);
  assign s_24 = s_1671?s_25:s_1670;
  assign s_25 = s_26[53:1];
  assign s_26 = s_1657?s_27:s_1656;
  dq #(54, 1) dq_s_27 (clk, s_27, s_28);
  assign s_28 = s_29 + s_1655;
  assign s_29 = s_30;
  assign s_30 = s_31[105:53];
  dq #(106, 1) dq_s_31 (clk, s_31, s_32);
  assign s_32 = s_33 << s_204;
  dq #(106, 2) dq_s_33 (clk, s_33, s_34);
  dq #(106, 1) dq_s_34 (clk, s_34, s_35);
  assign s_35 = s_36 >> s_189;
  assign s_36 = s_37[105:0];
  assign s_37 = {s_38,s_172};
  assign s_38 = s_39[16:0];
  dq #(49, 1) dq_s_39 (clk, s_39, s_40);
  assign s_40 = s_41;
  assign s_41 = s_42 + s_69;
  dq #(34, 14) dq_s_42 (clk, s_42, s_43);
  assign s_43 = s_44 * s_57;
  assign s_44 = s_45;
  assign s_45 = s_46[67:51];
  assign s_46 = s_47;
  assign s_47 = {s_48,s_56};
  assign s_48 = s_51?s_49:s_50;
  assign s_49 = 1'd0;
  assign s_50 = 1'd1;
  assign s_51 = s_52 == s_55;
  assign s_52 = s_53 - s_54;
  assign s_53 = s_5[62:52];
  assign s_54 = 10'd1023;
  assign s_55 = -11'd1023;
  assign s_56 = s_5[51:0];
  assign s_57 = s_58[67:51];
  assign s_58 = s_59;
  assign s_59 = {s_60,s_68};
  assign s_60 = s_63?s_61:s_62;
  assign s_61 = 1'd0;
  assign s_62 = 1'd1;
  assign s_63 = s_64 == s_67;
  assign s_64 = s_65 - s_66;
  assign s_65 = s_7[62:52];
  assign s_66 = 10'd1023;
  assign s_67 = -11'd1023;
  assign s_68 = s_7[51:0];
  assign s_69 = s_70 >> s_171;
  dq #(48, 1) dq_s_70 (clk, s_70, s_71);
  assign s_71 = s_72;
  assign s_72 = s_73 + s_77;
  dq #(34, 13) dq_s_73 (clk, s_73, s_74);
  assign s_74 = s_75 * s_76;
  assign s_75 = s_45;
  assign s_76 = s_58[50:34];
  dq #(47, 1) dq_s_77 (clk, s_77, s_78);
  assign s_78 = s_79;
  assign s_79 = s_80 + s_84;
  dq #(34, 12) dq_s_80 (clk, s_80, s_81);
  assign s_81 = s_82 * s_57;
  assign s_82 = s_83;
  assign s_83 = s_46[50:34];
  assign s_84 = s_85 >> s_170;
  dq #(46, 1) dq_s_85 (clk, s_85, s_86);
  assign s_86 = s_87;
  assign s_87 = s_88 + s_92;
  dq #(34, 11) dq_s_88 (clk, s_88, s_89);
  assign s_89 = s_90 * s_91;
  assign s_90 = s_45;
  assign s_91 = s_58[33:17];
  dq #(45, 1) dq_s_92 (clk, s_92, s_93);
  assign s_93 = s_94;
  assign s_94 = s_95 + s_98;
  dq #(34, 10) dq_s_95 (clk, s_95, s_96);
  assign s_96 = s_97 * s_76;
  assign s_97 = s_83;
  dq #(44, 1) dq_s_98 (clk, s_98, s_99);
  assign s_99 = s_100;
  assign s_100 = s_101 + s_105;
  dq #(34, 9) dq_s_101 (clk, s_101, s_102);
  assign s_102 = s_103 * s_57;
  assign s_103 = s_104;
  assign s_104 = s_46[33:17];
  assign s_105 = s_106 >> s_169;
  dq #(43, 1) dq_s_106 (clk, s_106, s_107);
  assign s_107 = s_108;
  assign s_108 = s_109 + s_113;
  dq #(34, 8) dq_s_109 (clk, s_109, s_110);
  assign s_110 = s_111 * s_112;
  assign s_111 = s_45;
  assign s_112 = s_58[16:0];
  dq #(42, 1) dq_s_113 (clk, s_113, s_114);
  assign s_114 = s_115;
  assign s_115 = s_116 + s_119;
  dq #(34, 7) dq_s_116 (clk, s_116, s_117);
  assign s_117 = s_118 * s_91;
  assign s_118 = s_83;
  dq #(41, 1) dq_s_119 (clk, s_119, s_120);
  assign s_120 = s_121;
  assign s_121 = s_122 + s_125;
  dq #(34, 6) dq_s_122 (clk, s_122, s_123);
  assign s_123 = s_124 * s_76;
  assign s_124 = s_104;
  dq #(40, 1) dq_s_125 (clk, s_125, s_126);
  assign s_126 = s_127;
  assign s_127 = s_128 + s_132;
  dq #(34, 5) dq_s_128 (clk, s_128, s_129);
  assign s_129 = s_130 * s_57;
  assign s_130 = s_131;
  assign s_131 = s_46[16:0];
  assign s_132 = s_133 >> s_168;
  dq #(39, 1) dq_s_133 (clk, s_133, s_134);
  assign s_134 = s_135;
  assign s_135 = s_136 + s_139;
  dq #(34, 4) dq_s_136 (clk, s_136, s_137);
  assign s_137 = s_138 * s_112;
  assign s_138 = s_83;
  dq #(38, 1) dq_s_139 (clk, s_139, s_140);
  assign s_140 = s_141;
  assign s_141 = s_142 + s_145;
  dq #(34, 3) dq_s_142 (clk, s_142, s_143);
  assign s_143 = s_144 * s_91;
  assign s_144 = s_104;
  dq #(37, 1) dq_s_145 (clk, s_145, s_146);
  assign s_146 = s_147;
  assign s_147 = s_148 + s_151;
  dq #(34, 2) dq_s_148 (clk, s_148, s_149);
  assign s_149 = s_150 * s_76;
  assign s_150 = s_131;
  assign s_151 = s_152 >> s_167;
  dq #(36, 1) dq_s_152 (clk, s_152, s_153);
  assign s_153 = s_154;
  assign s_154 = s_155 + s_158;
  dq #(34, 1) dq_s_155 (clk, s_155, s_156);
  assign s_156 = s_157 * s_112;
  assign s_157 = s_104;
  dq #(35, 1) dq_s_158 (clk, s_158, s_159);
  assign s_159 = s_160;
  assign s_160 = s_161 + s_163;
  assign s_161 = s_162 * s_91;
  assign s_162 = s_131;
  assign s_163 = s_164 >> s_166;
  assign s_164 = s_165 * s_112;
  assign s_165 = s_131;
  assign s_166 = 5'd17;
  assign s_167 = 5'd17;
  assign s_168 = 5'd17;
  assign s_169 = 5'd17;
  assign s_170 = 5'd17;
  assign s_171 = 5'd17;
  dq #(102, 1) dq_s_172 (clk, s_172, s_173);
  assign s_173 = {s_174,s_175};
  assign s_174 = s_70[16:0];
  dq #(85, 2) dq_s_175 (clk, s_175, s_176);
  assign s_176 = {s_177,s_178};
  assign s_177 = s_85[16:0];
  dq #(68, 3) dq_s_178 (clk, s_178, s_179);
  assign s_179 = {s_180,s_181};
  assign s_180 = s_106[16:0];
  dq #(51, 4) dq_s_181 (clk, s_181, s_182);
  assign s_182 = {s_183,s_184};
  assign s_183 = s_133[16:0];
  dq #(34, 3) dq_s_184 (clk, s_184, s_185);
  assign s_185 = {s_186,s_187};
  assign s_186 = s_152[16:0];
  dq #(17, 2) dq_s_187 (clk, s_187, s_188);
  assign s_188 = s_164[16:0];
  dq #(13, 15) dq_s_189 (clk, s_189, s_190);
  assign s_190 = s_203?s_191:s_192;
  assign s_191 = 1'd0;
  assign s_192 = s_193 - s_194;
  assign s_193 = -13'd1022;
  assign s_194 = s_195 + s_202;
  assign s_195 = s_196 + s_199;
  assign s_196 = $signed(s_197);
  assign s_197 = s_51?s_198:s_52;
  assign s_198 = -11'd1022;
  assign s_199 = $signed(s_200);
  assign s_200 = s_63?s_201:s_64;
  assign s_201 = -11'd1022;
  assign s_202 = 1'd1;
  assign s_203 = s_192[12];
  dq #(13, 1) dq_s_204 (clk, s_204, s_205);
  assign s_205 = s_1652?s_206:s_1647;
  dq #(8, 1) dq_s_206 (clk, s_206, s_207);
  assign s_207 = {s_208,s_1641};
  assign s_208 = s_209 & s_947;
  assign s_209 = s_210[6];
  assign s_210 = {s_211,s_941};
  assign s_211 = s_212 & s_599;
  assign s_212 = s_213[5];
  assign s_213 = {s_214,s_593};
  assign s_214 = s_215 & s_427;
  assign s_215 = s_216[4];
  assign s_216 = {s_217,s_421};
  assign s_217 = s_218 & s_343;
  assign s_218 = s_219[3];
  assign s_219 = {s_220,s_337};
  assign s_220 = s_221 & s_303;
  assign s_221 = s_222[2];
  assign s_222 = {s_223,s_297};
  assign s_223 = s_224 & s_285;
  assign s_224 = s_225[1];
  assign s_225 = {s_226,s_281};
  assign s_226 = s_227 & s_279;
  assign s_227 = ~s_228;
  assign s_228 = s_229[1];
  assign s_229 = s_230[3:2];
  assign s_230 = s_231[7:4];
  assign s_231 = s_232[15:8];
  assign s_232 = s_233[31:16];
  assign s_233 = s_234[63:32];
  assign s_234 = s_235[127:64];
  assign s_235 = {s_236,s_278};
  assign s_236 = {s_237,s_277};
  assign s_237 = {s_238,s_276};
  assign s_238 = {s_239,s_275};
  assign s_239 = {s_240,s_274};
  assign s_240 = {s_241,s_273};
  assign s_241 = {s_242,s_272};
  assign s_242 = {s_243,s_271};
  assign s_243 = {s_244,s_270};
  assign s_244 = {s_245,s_269};
  assign s_245 = {s_246,s_268};
  assign s_246 = {s_247,s_267};
  assign s_247 = {s_248,s_266};
  assign s_248 = {s_249,s_265};
  assign s_249 = {s_250,s_264};
  assign s_250 = {s_251,s_263};
  assign s_251 = {s_252,s_262};
  assign s_252 = {s_253,s_261};
  assign s_253 = {s_254,s_260};
  assign s_254 = {s_255,s_259};
  assign s_255 = {s_256,s_258};
  assign s_256 = {s_34,s_257};
  assign s_257 = 1'd1;
  assign s_258 = 1'd1;
  assign s_259 = 1'd1;
  assign s_260 = 1'd1;
  assign s_261 = 1'd1;
  assign s_262 = 1'd1;
  assign s_263 = 1'd1;
  assign s_264 = 1'd1;
  assign s_265 = 1'd1;
  assign s_266 = 1'd1;
  assign s_267 = 1'd1;
  assign s_268 = 1'd1;
  assign s_269 = 1'd1;
  assign s_270 = 1'd1;
  assign s_271 = 1'd1;
  assign s_272 = 1'd1;
  assign s_273 = 1'd1;
  assign s_274 = 1'd1;
  assign s_275 = 1'd1;
  assign s_276 = 1'd1;
  assign s_277 = 1'd1;
  assign s_278 = 1'd1;
  assign s_279 = ~s_280;
  assign s_280 = s_229[0];
  assign s_281 = s_282 & s_284;
  assign s_282 = ~s_283;
  assign s_283 = s_229[1];
  assign s_284 = s_229[0];
  assign s_285 = s_286[1];
  assign s_286 = {s_287,s_293};
  assign s_287 = s_288 & s_291;
  assign s_288 = ~s_289;
  assign s_289 = s_290[1];
  assign s_290 = s_230[1:0];
  assign s_291 = ~s_292;
  assign s_292 = s_290[0];
  assign s_293 = s_294 & s_296;
  assign s_294 = ~s_295;
  assign s_295 = s_290[1];
  assign s_296 = s_290[0];
  assign s_297 = {s_298,s_300};
  assign s_298 = s_224 & s_299;
  assign s_299 = ~s_285;
  assign s_300 = s_224?s_301:s_302;
  assign s_301 = s_286[0:0];
  assign s_302 = s_225[0:0];
  assign s_303 = s_304[2];
  assign s_304 = {s_305,s_331};
  assign s_305 = s_306 & s_319;
  assign s_306 = s_307[1];
  assign s_307 = {s_308,s_315};
  assign s_308 = s_309 & s_313;
  assign s_309 = ~s_310;
  assign s_310 = s_311[1];
  assign s_311 = s_312[3:2];
  assign s_312 = s_231[3:0];
  assign s_313 = ~s_314;
  assign s_314 = s_311[0];
  assign s_315 = s_316 & s_318;
  assign s_316 = ~s_317;
  assign s_317 = s_311[1];
  assign s_318 = s_311[0];
  assign s_319 = s_320[1];
  assign s_320 = {s_321,s_327};
  assign s_321 = s_322 & s_325;
  assign s_322 = ~s_323;
  assign s_323 = s_324[1];
  assign s_324 = s_312[1:0];
  assign s_325 = ~s_326;
  assign s_326 = s_324[0];
  assign s_327 = s_328 & s_330;
  assign s_328 = ~s_329;
  assign s_329 = s_324[1];
  assign s_330 = s_324[0];
  assign s_331 = {s_332,s_334};
  assign s_332 = s_306 & s_333;
  assign s_333 = ~s_319;
  assign s_334 = s_306?s_335:s_336;
  assign s_335 = s_320[0:0];
  assign s_336 = s_307[0:0];
  assign s_337 = {s_338,s_340};
  assign s_338 = s_221 & s_339;
  assign s_339 = ~s_303;
  assign s_340 = s_221?s_341:s_342;
  assign s_341 = s_304[1:0];
  assign s_342 = s_222[1:0];
  assign s_343 = s_344[3];
  assign s_344 = {s_345,s_415};
  assign s_345 = s_346 & s_381;
  assign s_346 = s_347[2];
  assign s_347 = {s_348,s_375};
  assign s_348 = s_349 & s_363;
  assign s_349 = s_350[1];
  assign s_350 = {s_351,s_359};
  assign s_351 = s_352 & s_357;
  assign s_352 = ~s_353;
  assign s_353 = s_354[1];
  assign s_354 = s_355[3:2];
  assign s_355 = s_356[7:4];
  assign s_356 = s_232[7:0];
  assign s_357 = ~s_358;
  assign s_358 = s_354[0];
  assign s_359 = s_360 & s_362;
  assign s_360 = ~s_361;
  assign s_361 = s_354[1];
  assign s_362 = s_354[0];
  assign s_363 = s_364[1];
  assign s_364 = {s_365,s_371};
  assign s_365 = s_366 & s_369;
  assign s_366 = ~s_367;
  assign s_367 = s_368[1];
  assign s_368 = s_355[1:0];
  assign s_369 = ~s_370;
  assign s_370 = s_368[0];
  assign s_371 = s_372 & s_374;
  assign s_372 = ~s_373;
  assign s_373 = s_368[1];
  assign s_374 = s_368[0];
  assign s_375 = {s_376,s_378};
  assign s_376 = s_349 & s_377;
  assign s_377 = ~s_363;
  assign s_378 = s_349?s_379:s_380;
  assign s_379 = s_364[0:0];
  assign s_380 = s_350[0:0];
  assign s_381 = s_382[2];
  assign s_382 = {s_383,s_409};
  assign s_383 = s_384 & s_397;
  assign s_384 = s_385[1];
  assign s_385 = {s_386,s_393};
  assign s_386 = s_387 & s_391;
  assign s_387 = ~s_388;
  assign s_388 = s_389[1];
  assign s_389 = s_390[3:2];
  assign s_390 = s_356[3:0];
  assign s_391 = ~s_392;
  assign s_392 = s_389[0];
  assign s_393 = s_394 & s_396;
  assign s_394 = ~s_395;
  assign s_395 = s_389[1];
  assign s_396 = s_389[0];
  assign s_397 = s_398[1];
  assign s_398 = {s_399,s_405};
  assign s_399 = s_400 & s_403;
  assign s_400 = ~s_401;
  assign s_401 = s_402[1];
  assign s_402 = s_390[1:0];
  assign s_403 = ~s_404;
  assign s_404 = s_402[0];
  assign s_405 = s_406 & s_408;
  assign s_406 = ~s_407;
  assign s_407 = s_402[1];
  assign s_408 = s_402[0];
  assign s_409 = {s_410,s_412};
  assign s_410 = s_384 & s_411;
  assign s_411 = ~s_397;
  assign s_412 = s_384?s_413:s_414;
  assign s_413 = s_398[0:0];
  assign s_414 = s_385[0:0];
  assign s_415 = {s_416,s_418};
  assign s_416 = s_346 & s_417;
  assign s_417 = ~s_381;
  assign s_418 = s_346?s_419:s_420;
  assign s_419 = s_382[1:0];
  assign s_420 = s_347[1:0];
  assign s_421 = {s_422,s_424};
  assign s_422 = s_218 & s_423;
  assign s_423 = ~s_343;
  assign s_424 = s_218?s_425:s_426;
  assign s_425 = s_344[2:0];
  assign s_426 = s_219[2:0];
  assign s_427 = s_428[4];
  assign s_428 = {s_429,s_587};
  assign s_429 = s_430 & s_509;
  assign s_430 = s_431[3];
  assign s_431 = {s_432,s_503};
  assign s_432 = s_433 & s_469;
  assign s_433 = s_434[2];
  assign s_434 = {s_435,s_463};
  assign s_435 = s_436 & s_451;
  assign s_436 = s_437[1];
  assign s_437 = {s_438,s_447};
  assign s_438 = s_439 & s_445;
  assign s_439 = ~s_440;
  assign s_440 = s_441[1];
  assign s_441 = s_442[3:2];
  assign s_442 = s_443[7:4];
  assign s_443 = s_444[15:8];
  assign s_444 = s_233[15:0];
  assign s_445 = ~s_446;
  assign s_446 = s_441[0];
  assign s_447 = s_448 & s_450;
  assign s_448 = ~s_449;
  assign s_449 = s_441[1];
  assign s_450 = s_441[0];
  assign s_451 = s_452[1];
  assign s_452 = {s_453,s_459};
  assign s_453 = s_454 & s_457;
  assign s_454 = ~s_455;
  assign s_455 = s_456[1];
  assign s_456 = s_442[1:0];
  assign s_457 = ~s_458;
  assign s_458 = s_456[0];
  assign s_459 = s_460 & s_462;
  assign s_460 = ~s_461;
  assign s_461 = s_456[1];
  assign s_462 = s_456[0];
  assign s_463 = {s_464,s_466};
  assign s_464 = s_436 & s_465;
  assign s_465 = ~s_451;
  assign s_466 = s_436?s_467:s_468;
  assign s_467 = s_452[0:0];
  assign s_468 = s_437[0:0];
  assign s_469 = s_470[2];
  assign s_470 = {s_471,s_497};
  assign s_471 = s_472 & s_485;
  assign s_472 = s_473[1];
  assign s_473 = {s_474,s_481};
  assign s_474 = s_475 & s_479;
  assign s_475 = ~s_476;
  assign s_476 = s_477[1];
  assign s_477 = s_478[3:2];
  assign s_478 = s_443[3:0];
  assign s_479 = ~s_480;
  assign s_480 = s_477[0];
  assign s_481 = s_482 & s_484;
  assign s_482 = ~s_483;
  assign s_483 = s_477[1];
  assign s_484 = s_477[0];
  assign s_485 = s_486[1];
  assign s_486 = {s_487,s_493};
  assign s_487 = s_488 & s_491;
  assign s_488 = ~s_489;
  assign s_489 = s_490[1];
  assign s_490 = s_478[1:0];
  assign s_491 = ~s_492;
  assign s_492 = s_490[0];
  assign s_493 = s_494 & s_496;
  assign s_494 = ~s_495;
  assign s_495 = s_490[1];
  assign s_496 = s_490[0];
  assign s_497 = {s_498,s_500};
  assign s_498 = s_472 & s_499;
  assign s_499 = ~s_485;
  assign s_500 = s_472?s_501:s_502;
  assign s_501 = s_486[0:0];
  assign s_502 = s_473[0:0];
  assign s_503 = {s_504,s_506};
  assign s_504 = s_433 & s_505;
  assign s_505 = ~s_469;
  assign s_506 = s_433?s_507:s_508;
  assign s_507 = s_470[1:0];
  assign s_508 = s_434[1:0];
  assign s_509 = s_510[3];
  assign s_510 = {s_511,s_581};
  assign s_511 = s_512 & s_547;
  assign s_512 = s_513[2];
  assign s_513 = {s_514,s_541};
  assign s_514 = s_515 & s_529;
  assign s_515 = s_516[1];
  assign s_516 = {s_517,s_525};
  assign s_517 = s_518 & s_523;
  assign s_518 = ~s_519;
  assign s_519 = s_520[1];
  assign s_520 = s_521[3:2];
  assign s_521 = s_522[7:4];
  assign s_522 = s_444[7:0];
  assign s_523 = ~s_524;
  assign s_524 = s_520[0];
  assign s_525 = s_526 & s_528;
  assign s_526 = ~s_527;
  assign s_527 = s_520[1];
  assign s_528 = s_520[0];
  assign s_529 = s_530[1];
  assign s_530 = {s_531,s_537};
  assign s_531 = s_532 & s_535;
  assign s_532 = ~s_533;
  assign s_533 = s_534[1];
  assign s_534 = s_521[1:0];
  assign s_535 = ~s_536;
  assign s_536 = s_534[0];
  assign s_537 = s_538 & s_540;
  assign s_538 = ~s_539;
  assign s_539 = s_534[1];
  assign s_540 = s_534[0];
  assign s_541 = {s_542,s_544};
  assign s_542 = s_515 & s_543;
  assign s_543 = ~s_529;
  assign s_544 = s_515?s_545:s_546;
  assign s_545 = s_530[0:0];
  assign s_546 = s_516[0:0];
  assign s_547 = s_548[2];
  assign s_548 = {s_549,s_575};
  assign s_549 = s_550 & s_563;
  assign s_550 = s_551[1];
  assign s_551 = {s_552,s_559};
  assign s_552 = s_553 & s_557;
  assign s_553 = ~s_554;
  assign s_554 = s_555[1];
  assign s_555 = s_556[3:2];
  assign s_556 = s_522[3:0];
  assign s_557 = ~s_558;
  assign s_558 = s_555[0];
  assign s_559 = s_560 & s_562;
  assign s_560 = ~s_561;
  assign s_561 = s_555[1];
  assign s_562 = s_555[0];
  assign s_563 = s_564[1];
  assign s_564 = {s_565,s_571};
  assign s_565 = s_566 & s_569;
  assign s_566 = ~s_567;
  assign s_567 = s_568[1];
  assign s_568 = s_556[1:0];
  assign s_569 = ~s_570;
  assign s_570 = s_568[0];
  assign s_571 = s_572 & s_574;
  assign s_572 = ~s_573;
  assign s_573 = s_568[1];
  assign s_574 = s_568[0];
  assign s_575 = {s_576,s_578};
  assign s_576 = s_550 & s_577;
  assign s_577 = ~s_563;
  assign s_578 = s_550?s_579:s_580;
  assign s_579 = s_564[0:0];
  assign s_580 = s_551[0:0];
  assign s_581 = {s_582,s_584};
  assign s_582 = s_512 & s_583;
  assign s_583 = ~s_547;
  assign s_584 = s_512?s_585:s_586;
  assign s_585 = s_548[1:0];
  assign s_586 = s_513[1:0];
  assign s_587 = {s_588,s_590};
  assign s_588 = s_430 & s_589;
  assign s_589 = ~s_509;
  assign s_590 = s_430?s_591:s_592;
  assign s_591 = s_510[2:0];
  assign s_592 = s_431[2:0];
  assign s_593 = {s_594,s_596};
  assign s_594 = s_215 & s_595;
  assign s_595 = ~s_427;
  assign s_596 = s_215?s_597:s_598;
  assign s_597 = s_428[3:0];
  assign s_598 = s_216[3:0];
  assign s_599 = s_600[5];
  assign s_600 = {s_601,s_935};
  assign s_601 = s_602 & s_769;
  assign s_602 = s_603[4];
  assign s_603 = {s_604,s_763};
  assign s_604 = s_605 & s_685;
  assign s_605 = s_606[3];
  assign s_606 = {s_607,s_679};
  assign s_607 = s_608 & s_645;
  assign s_608 = s_609[2];
  assign s_609 = {s_610,s_639};
  assign s_610 = s_611 & s_627;
  assign s_611 = s_612[1];
  assign s_612 = {s_613,s_623};
  assign s_613 = s_614 & s_621;
  assign s_614 = ~s_615;
  assign s_615 = s_616[1];
  assign s_616 = s_617[3:2];
  assign s_617 = s_618[7:4];
  assign s_618 = s_619[15:8];
  assign s_619 = s_620[31:16];
  assign s_620 = s_234[31:0];
  assign s_621 = ~s_622;
  assign s_622 = s_616[0];
  assign s_623 = s_624 & s_626;
  assign s_624 = ~s_625;
  assign s_625 = s_616[1];
  assign s_626 = s_616[0];
  assign s_627 = s_628[1];
  assign s_628 = {s_629,s_635};
  assign s_629 = s_630 & s_633;
  assign s_630 = ~s_631;
  assign s_631 = s_632[1];
  assign s_632 = s_617[1:0];
  assign s_633 = ~s_634;
  assign s_634 = s_632[0];
  assign s_635 = s_636 & s_638;
  assign s_636 = ~s_637;
  assign s_637 = s_632[1];
  assign s_638 = s_632[0];
  assign s_639 = {s_640,s_642};
  assign s_640 = s_611 & s_641;
  assign s_641 = ~s_627;
  assign s_642 = s_611?s_643:s_644;
  assign s_643 = s_628[0:0];
  assign s_644 = s_612[0:0];
  assign s_645 = s_646[2];
  assign s_646 = {s_647,s_673};
  assign s_647 = s_648 & s_661;
  assign s_648 = s_649[1];
  assign s_649 = {s_650,s_657};
  assign s_650 = s_651 & s_655;
  assign s_651 = ~s_652;
  assign s_652 = s_653[1];
  assign s_653 = s_654[3:2];
  assign s_654 = s_618[3:0];
  assign s_655 = ~s_656;
  assign s_656 = s_653[0];
  assign s_657 = s_658 & s_660;
  assign s_658 = ~s_659;
  assign s_659 = s_653[1];
  assign s_660 = s_653[0];
  assign s_661 = s_662[1];
  assign s_662 = {s_663,s_669};
  assign s_663 = s_664 & s_667;
  assign s_664 = ~s_665;
  assign s_665 = s_666[1];
  assign s_666 = s_654[1:0];
  assign s_667 = ~s_668;
  assign s_668 = s_666[0];
  assign s_669 = s_670 & s_672;
  assign s_670 = ~s_671;
  assign s_671 = s_666[1];
  assign s_672 = s_666[0];
  assign s_673 = {s_674,s_676};
  assign s_674 = s_648 & s_675;
  assign s_675 = ~s_661;
  assign s_676 = s_648?s_677:s_678;
  assign s_677 = s_662[0:0];
  assign s_678 = s_649[0:0];
  assign s_679 = {s_680,s_682};
  assign s_680 = s_608 & s_681;
  assign s_681 = ~s_645;
  assign s_682 = s_608?s_683:s_684;
  assign s_683 = s_646[1:0];
  assign s_684 = s_609[1:0];
  assign s_685 = s_686[3];
  assign s_686 = {s_687,s_757};
  assign s_687 = s_688 & s_723;
  assign s_688 = s_689[2];
  assign s_689 = {s_690,s_717};
  assign s_690 = s_691 & s_705;
  assign s_691 = s_692[1];
  assign s_692 = {s_693,s_701};
  assign s_693 = s_694 & s_699;
  assign s_694 = ~s_695;
  assign s_695 = s_696[1];
  assign s_696 = s_697[3:2];
  assign s_697 = s_698[7:4];
  assign s_698 = s_619[7:0];
  assign s_699 = ~s_700;
  assign s_700 = s_696[0];
  assign s_701 = s_702 & s_704;
  assign s_702 = ~s_703;
  assign s_703 = s_696[1];
  assign s_704 = s_696[0];
  assign s_705 = s_706[1];
  assign s_706 = {s_707,s_713};
  assign s_707 = s_708 & s_711;
  assign s_708 = ~s_709;
  assign s_709 = s_710[1];
  assign s_710 = s_697[1:0];
  assign s_711 = ~s_712;
  assign s_712 = s_710[0];
  assign s_713 = s_714 & s_716;
  assign s_714 = ~s_715;
  assign s_715 = s_710[1];
  assign s_716 = s_710[0];
  assign s_717 = {s_718,s_720};
  assign s_718 = s_691 & s_719;
  assign s_719 = ~s_705;
  assign s_720 = s_691?s_721:s_722;
  assign s_721 = s_706[0:0];
  assign s_722 = s_692[0:0];
  assign s_723 = s_724[2];
  assign s_724 = {s_725,s_751};
  assign s_725 = s_726 & s_739;
  assign s_726 = s_727[1];
  assign s_727 = {s_728,s_735};
  assign s_728 = s_729 & s_733;
  assign s_729 = ~s_730;
  assign s_730 = s_731[1];
  assign s_731 = s_732[3:2];
  assign s_732 = s_698[3:0];
  assign s_733 = ~s_734;
  assign s_734 = s_731[0];
  assign s_735 = s_736 & s_738;
  assign s_736 = ~s_737;
  assign s_737 = s_731[1];
  assign s_738 = s_731[0];
  assign s_739 = s_740[1];
  assign s_740 = {s_741,s_747};
  assign s_741 = s_742 & s_745;
  assign s_742 = ~s_743;
  assign s_743 = s_744[1];
  assign s_744 = s_732[1:0];
  assign s_745 = ~s_746;
  assign s_746 = s_744[0];
  assign s_747 = s_748 & s_750;
  assign s_748 = ~s_749;
  assign s_749 = s_744[1];
  assign s_750 = s_744[0];
  assign s_751 = {s_752,s_754};
  assign s_752 = s_726 & s_753;
  assign s_753 = ~s_739;
  assign s_754 = s_726?s_755:s_756;
  assign s_755 = s_740[0:0];
  assign s_756 = s_727[0:0];
  assign s_757 = {s_758,s_760};
  assign s_758 = s_688 & s_759;
  assign s_759 = ~s_723;
  assign s_760 = s_688?s_761:s_762;
  assign s_761 = s_724[1:0];
  assign s_762 = s_689[1:0];
  assign s_763 = {s_764,s_766};
  assign s_764 = s_605 & s_765;
  assign s_765 = ~s_685;
  assign s_766 = s_605?s_767:s_768;
  assign s_767 = s_686[2:0];
  assign s_768 = s_606[2:0];
  assign s_769 = s_770[4];
  assign s_770 = {s_771,s_929};
  assign s_771 = s_772 & s_851;
  assign s_772 = s_773[3];
  assign s_773 = {s_774,s_845};
  assign s_774 = s_775 & s_811;
  assign s_775 = s_776[2];
  assign s_776 = {s_777,s_805};
  assign s_777 = s_778 & s_793;
  assign s_778 = s_779[1];
  assign s_779 = {s_780,s_789};
  assign s_780 = s_781 & s_787;
  assign s_781 = ~s_782;
  assign s_782 = s_783[1];
  assign s_783 = s_784[3:2];
  assign s_784 = s_785[7:4];
  assign s_785 = s_786[15:8];
  assign s_786 = s_620[15:0];
  assign s_787 = ~s_788;
  assign s_788 = s_783[0];
  assign s_789 = s_790 & s_792;
  assign s_790 = ~s_791;
  assign s_791 = s_783[1];
  assign s_792 = s_783[0];
  assign s_793 = s_794[1];
  assign s_794 = {s_795,s_801};
  assign s_795 = s_796 & s_799;
  assign s_796 = ~s_797;
  assign s_797 = s_798[1];
  assign s_798 = s_784[1:0];
  assign s_799 = ~s_800;
  assign s_800 = s_798[0];
  assign s_801 = s_802 & s_804;
  assign s_802 = ~s_803;
  assign s_803 = s_798[1];
  assign s_804 = s_798[0];
  assign s_805 = {s_806,s_808};
  assign s_806 = s_778 & s_807;
  assign s_807 = ~s_793;
  assign s_808 = s_778?s_809:s_810;
  assign s_809 = s_794[0:0];
  assign s_810 = s_779[0:0];
  assign s_811 = s_812[2];
  assign s_812 = {s_813,s_839};
  assign s_813 = s_814 & s_827;
  assign s_814 = s_815[1];
  assign s_815 = {s_816,s_823};
  assign s_816 = s_817 & s_821;
  assign s_817 = ~s_818;
  assign s_818 = s_819[1];
  assign s_819 = s_820[3:2];
  assign s_820 = s_785[3:0];
  assign s_821 = ~s_822;
  assign s_822 = s_819[0];
  assign s_823 = s_824 & s_826;
  assign s_824 = ~s_825;
  assign s_825 = s_819[1];
  assign s_826 = s_819[0];
  assign s_827 = s_828[1];
  assign s_828 = {s_829,s_835};
  assign s_829 = s_830 & s_833;
  assign s_830 = ~s_831;
  assign s_831 = s_832[1];
  assign s_832 = s_820[1:0];
  assign s_833 = ~s_834;
  assign s_834 = s_832[0];
  assign s_835 = s_836 & s_838;
  assign s_836 = ~s_837;
  assign s_837 = s_832[1];
  assign s_838 = s_832[0];
  assign s_839 = {s_840,s_842};
  assign s_840 = s_814 & s_841;
  assign s_841 = ~s_827;
  assign s_842 = s_814?s_843:s_844;
  assign s_843 = s_828[0:0];
  assign s_844 = s_815[0:0];
  assign s_845 = {s_846,s_848};
  assign s_846 = s_775 & s_847;
  assign s_847 = ~s_811;
  assign s_848 = s_775?s_849:s_850;
  assign s_849 = s_812[1:0];
  assign s_850 = s_776[1:0];
  assign s_851 = s_852[3];
  assign s_852 = {s_853,s_923};
  assign s_853 = s_854 & s_889;
  assign s_854 = s_855[2];
  assign s_855 = {s_856,s_883};
  assign s_856 = s_857 & s_871;
  assign s_857 = s_858[1];
  assign s_858 = {s_859,s_867};
  assign s_859 = s_860 & s_865;
  assign s_860 = ~s_861;
  assign s_861 = s_862[1];
  assign s_862 = s_863[3:2];
  assign s_863 = s_864[7:4];
  assign s_864 = s_786[7:0];
  assign s_865 = ~s_866;
  assign s_866 = s_862[0];
  assign s_867 = s_868 & s_870;
  assign s_868 = ~s_869;
  assign s_869 = s_862[1];
  assign s_870 = s_862[0];
  assign s_871 = s_872[1];
  assign s_872 = {s_873,s_879};
  assign s_873 = s_874 & s_877;
  assign s_874 = ~s_875;
  assign s_875 = s_876[1];
  assign s_876 = s_863[1:0];
  assign s_877 = ~s_878;
  assign s_878 = s_876[0];
  assign s_879 = s_880 & s_882;
  assign s_880 = ~s_881;
  assign s_881 = s_876[1];
  assign s_882 = s_876[0];
  assign s_883 = {s_884,s_886};
  assign s_884 = s_857 & s_885;
  assign s_885 = ~s_871;
  assign s_886 = s_857?s_887:s_888;
  assign s_887 = s_872[0:0];
  assign s_888 = s_858[0:0];
  assign s_889 = s_890[2];
  assign s_890 = {s_891,s_917};
  assign s_891 = s_892 & s_905;
  assign s_892 = s_893[1];
  assign s_893 = {s_894,s_901};
  assign s_894 = s_895 & s_899;
  assign s_895 = ~s_896;
  assign s_896 = s_897[1];
  assign s_897 = s_898[3:2];
  assign s_898 = s_864[3:0];
  assign s_899 = ~s_900;
  assign s_900 = s_897[0];
  assign s_901 = s_902 & s_904;
  assign s_902 = ~s_903;
  assign s_903 = s_897[1];
  assign s_904 = s_897[0];
  assign s_905 = s_906[1];
  assign s_906 = {s_907,s_913};
  assign s_907 = s_908 & s_911;
  assign s_908 = ~s_909;
  assign s_909 = s_910[1];
  assign s_910 = s_898[1:0];
  assign s_911 = ~s_912;
  assign s_912 = s_910[0];
  assign s_913 = s_914 & s_916;
  assign s_914 = ~s_915;
  assign s_915 = s_910[1];
  assign s_916 = s_910[0];
  assign s_917 = {s_918,s_920};
  assign s_918 = s_892 & s_919;
  assign s_919 = ~s_905;
  assign s_920 = s_892?s_921:s_922;
  assign s_921 = s_906[0:0];
  assign s_922 = s_893[0:0];
  assign s_923 = {s_924,s_926};
  assign s_924 = s_854 & s_925;
  assign s_925 = ~s_889;
  assign s_926 = s_854?s_927:s_928;
  assign s_927 = s_890[1:0];
  assign s_928 = s_855[1:0];
  assign s_929 = {s_930,s_932};
  assign s_930 = s_772 & s_931;
  assign s_931 = ~s_851;
  assign s_932 = s_772?s_933:s_934;
  assign s_933 = s_852[2:0];
  assign s_934 = s_773[2:0];
  assign s_935 = {s_936,s_938};
  assign s_936 = s_602 & s_937;
  assign s_937 = ~s_769;
  assign s_938 = s_602?s_939:s_940;
  assign s_939 = s_770[3:0];
  assign s_940 = s_603[3:0];
  assign s_941 = {s_942,s_944};
  assign s_942 = s_212 & s_943;
  assign s_943 = ~s_599;
  assign s_944 = s_212?s_945:s_946;
  assign s_945 = s_600[4:0];
  assign s_946 = s_213[4:0];
  assign s_947 = s_948[6];
  assign s_948 = {s_949,s_1635};
  assign s_949 = s_950 & s_1293;
  assign s_950 = s_951[5];
  assign s_951 = {s_952,s_1287};
  assign s_952 = s_953 & s_1121;
  assign s_953 = s_954[4];
  assign s_954 = {s_955,s_1115};
  assign s_955 = s_956 & s_1037;
  assign s_956 = s_957[3];
  assign s_957 = {s_958,s_1031};
  assign s_958 = s_959 & s_997;
  assign s_959 = s_960[2];
  assign s_960 = {s_961,s_991};
  assign s_961 = s_962 & s_979;
  assign s_962 = s_963[1];
  assign s_963 = {s_964,s_975};
  assign s_964 = s_965 & s_973;
  assign s_965 = ~s_966;
  assign s_966 = s_967[1];
  assign s_967 = s_968[3:2];
  assign s_968 = s_969[7:4];
  assign s_969 = s_970[15:8];
  assign s_970 = s_971[31:16];
  assign s_971 = s_972[63:32];
  assign s_972 = s_235[63:0];
  assign s_973 = ~s_974;
  assign s_974 = s_967[0];
  assign s_975 = s_976 & s_978;
  assign s_976 = ~s_977;
  assign s_977 = s_967[1];
  assign s_978 = s_967[0];
  assign s_979 = s_980[1];
  assign s_980 = {s_981,s_987};
  assign s_981 = s_982 & s_985;
  assign s_982 = ~s_983;
  assign s_983 = s_984[1];
  assign s_984 = s_968[1:0];
  assign s_985 = ~s_986;
  assign s_986 = s_984[0];
  assign s_987 = s_988 & s_990;
  assign s_988 = ~s_989;
  assign s_989 = s_984[1];
  assign s_990 = s_984[0];
  assign s_991 = {s_992,s_994};
  assign s_992 = s_962 & s_993;
  assign s_993 = ~s_979;
  assign s_994 = s_962?s_995:s_996;
  assign s_995 = s_980[0:0];
  assign s_996 = s_963[0:0];
  assign s_997 = s_998[2];
  assign s_998 = {s_999,s_1025};
  assign s_999 = s_1000 & s_1013;
  assign s_1000 = s_1001[1];
  assign s_1001 = {s_1002,s_1009};
  assign s_1002 = s_1003 & s_1007;
  assign s_1003 = ~s_1004;
  assign s_1004 = s_1005[1];
  assign s_1005 = s_1006[3:2];
  assign s_1006 = s_969[3:0];
  assign s_1007 = ~s_1008;
  assign s_1008 = s_1005[0];
  assign s_1009 = s_1010 & s_1012;
  assign s_1010 = ~s_1011;
  assign s_1011 = s_1005[1];
  assign s_1012 = s_1005[0];
  assign s_1013 = s_1014[1];
  assign s_1014 = {s_1015,s_1021};
  assign s_1015 = s_1016 & s_1019;
  assign s_1016 = ~s_1017;
  assign s_1017 = s_1018[1];
  assign s_1018 = s_1006[1:0];
  assign s_1019 = ~s_1020;
  assign s_1020 = s_1018[0];
  assign s_1021 = s_1022 & s_1024;
  assign s_1022 = ~s_1023;
  assign s_1023 = s_1018[1];
  assign s_1024 = s_1018[0];
  assign s_1025 = {s_1026,s_1028};
  assign s_1026 = s_1000 & s_1027;
  assign s_1027 = ~s_1013;
  assign s_1028 = s_1000?s_1029:s_1030;
  assign s_1029 = s_1014[0:0];
  assign s_1030 = s_1001[0:0];
  assign s_1031 = {s_1032,s_1034};
  assign s_1032 = s_959 & s_1033;
  assign s_1033 = ~s_997;
  assign s_1034 = s_959?s_1035:s_1036;
  assign s_1035 = s_998[1:0];
  assign s_1036 = s_960[1:0];
  assign s_1037 = s_1038[3];
  assign s_1038 = {s_1039,s_1109};
  assign s_1039 = s_1040 & s_1075;
  assign s_1040 = s_1041[2];
  assign s_1041 = {s_1042,s_1069};
  assign s_1042 = s_1043 & s_1057;
  assign s_1043 = s_1044[1];
  assign s_1044 = {s_1045,s_1053};
  assign s_1045 = s_1046 & s_1051;
  assign s_1046 = ~s_1047;
  assign s_1047 = s_1048[1];
  assign s_1048 = s_1049[3:2];
  assign s_1049 = s_1050[7:4];
  assign s_1050 = s_970[7:0];
  assign s_1051 = ~s_1052;
  assign s_1052 = s_1048[0];
  assign s_1053 = s_1054 & s_1056;
  assign s_1054 = ~s_1055;
  assign s_1055 = s_1048[1];
  assign s_1056 = s_1048[0];
  assign s_1057 = s_1058[1];
  assign s_1058 = {s_1059,s_1065};
  assign s_1059 = s_1060 & s_1063;
  assign s_1060 = ~s_1061;
  assign s_1061 = s_1062[1];
  assign s_1062 = s_1049[1:0];
  assign s_1063 = ~s_1064;
  assign s_1064 = s_1062[0];
  assign s_1065 = s_1066 & s_1068;
  assign s_1066 = ~s_1067;
  assign s_1067 = s_1062[1];
  assign s_1068 = s_1062[0];
  assign s_1069 = {s_1070,s_1072};
  assign s_1070 = s_1043 & s_1071;
  assign s_1071 = ~s_1057;
  assign s_1072 = s_1043?s_1073:s_1074;
  assign s_1073 = s_1058[0:0];
  assign s_1074 = s_1044[0:0];
  assign s_1075 = s_1076[2];
  assign s_1076 = {s_1077,s_1103};
  assign s_1077 = s_1078 & s_1091;
  assign s_1078 = s_1079[1];
  assign s_1079 = {s_1080,s_1087};
  assign s_1080 = s_1081 & s_1085;
  assign s_1081 = ~s_1082;
  assign s_1082 = s_1083[1];
  assign s_1083 = s_1084[3:2];
  assign s_1084 = s_1050[3:0];
  assign s_1085 = ~s_1086;
  assign s_1086 = s_1083[0];
  assign s_1087 = s_1088 & s_1090;
  assign s_1088 = ~s_1089;
  assign s_1089 = s_1083[1];
  assign s_1090 = s_1083[0];
  assign s_1091 = s_1092[1];
  assign s_1092 = {s_1093,s_1099};
  assign s_1093 = s_1094 & s_1097;
  assign s_1094 = ~s_1095;
  assign s_1095 = s_1096[1];
  assign s_1096 = s_1084[1:0];
  assign s_1097 = ~s_1098;
  assign s_1098 = s_1096[0];
  assign s_1099 = s_1100 & s_1102;
  assign s_1100 = ~s_1101;
  assign s_1101 = s_1096[1];
  assign s_1102 = s_1096[0];
  assign s_1103 = {s_1104,s_1106};
  assign s_1104 = s_1078 & s_1105;
  assign s_1105 = ~s_1091;
  assign s_1106 = s_1078?s_1107:s_1108;
  assign s_1107 = s_1092[0:0];
  assign s_1108 = s_1079[0:0];
  assign s_1109 = {s_1110,s_1112};
  assign s_1110 = s_1040 & s_1111;
  assign s_1111 = ~s_1075;
  assign s_1112 = s_1040?s_1113:s_1114;
  assign s_1113 = s_1076[1:0];
  assign s_1114 = s_1041[1:0];
  assign s_1115 = {s_1116,s_1118};
  assign s_1116 = s_956 & s_1117;
  assign s_1117 = ~s_1037;
  assign s_1118 = s_956?s_1119:s_1120;
  assign s_1119 = s_1038[2:0];
  assign s_1120 = s_957[2:0];
  assign s_1121 = s_1122[4];
  assign s_1122 = {s_1123,s_1281};
  assign s_1123 = s_1124 & s_1203;
  assign s_1124 = s_1125[3];
  assign s_1125 = {s_1126,s_1197};
  assign s_1126 = s_1127 & s_1163;
  assign s_1127 = s_1128[2];
  assign s_1128 = {s_1129,s_1157};
  assign s_1129 = s_1130 & s_1145;
  assign s_1130 = s_1131[1];
  assign s_1131 = {s_1132,s_1141};
  assign s_1132 = s_1133 & s_1139;
  assign s_1133 = ~s_1134;
  assign s_1134 = s_1135[1];
  assign s_1135 = s_1136[3:2];
  assign s_1136 = s_1137[7:4];
  assign s_1137 = s_1138[15:8];
  assign s_1138 = s_971[15:0];
  assign s_1139 = ~s_1140;
  assign s_1140 = s_1135[0];
  assign s_1141 = s_1142 & s_1144;
  assign s_1142 = ~s_1143;
  assign s_1143 = s_1135[1];
  assign s_1144 = s_1135[0];
  assign s_1145 = s_1146[1];
  assign s_1146 = {s_1147,s_1153};
  assign s_1147 = s_1148 & s_1151;
  assign s_1148 = ~s_1149;
  assign s_1149 = s_1150[1];
  assign s_1150 = s_1136[1:0];
  assign s_1151 = ~s_1152;
  assign s_1152 = s_1150[0];
  assign s_1153 = s_1154 & s_1156;
  assign s_1154 = ~s_1155;
  assign s_1155 = s_1150[1];
  assign s_1156 = s_1150[0];
  assign s_1157 = {s_1158,s_1160};
  assign s_1158 = s_1130 & s_1159;
  assign s_1159 = ~s_1145;
  assign s_1160 = s_1130?s_1161:s_1162;
  assign s_1161 = s_1146[0:0];
  assign s_1162 = s_1131[0:0];
  assign s_1163 = s_1164[2];
  assign s_1164 = {s_1165,s_1191};
  assign s_1165 = s_1166 & s_1179;
  assign s_1166 = s_1167[1];
  assign s_1167 = {s_1168,s_1175};
  assign s_1168 = s_1169 & s_1173;
  assign s_1169 = ~s_1170;
  assign s_1170 = s_1171[1];
  assign s_1171 = s_1172[3:2];
  assign s_1172 = s_1137[3:0];
  assign s_1173 = ~s_1174;
  assign s_1174 = s_1171[0];
  assign s_1175 = s_1176 & s_1178;
  assign s_1176 = ~s_1177;
  assign s_1177 = s_1171[1];
  assign s_1178 = s_1171[0];
  assign s_1179 = s_1180[1];
  assign s_1180 = {s_1181,s_1187};
  assign s_1181 = s_1182 & s_1185;
  assign s_1182 = ~s_1183;
  assign s_1183 = s_1184[1];
  assign s_1184 = s_1172[1:0];
  assign s_1185 = ~s_1186;
  assign s_1186 = s_1184[0];
  assign s_1187 = s_1188 & s_1190;
  assign s_1188 = ~s_1189;
  assign s_1189 = s_1184[1];
  assign s_1190 = s_1184[0];
  assign s_1191 = {s_1192,s_1194};
  assign s_1192 = s_1166 & s_1193;
  assign s_1193 = ~s_1179;
  assign s_1194 = s_1166?s_1195:s_1196;
  assign s_1195 = s_1180[0:0];
  assign s_1196 = s_1167[0:0];
  assign s_1197 = {s_1198,s_1200};
  assign s_1198 = s_1127 & s_1199;
  assign s_1199 = ~s_1163;
  assign s_1200 = s_1127?s_1201:s_1202;
  assign s_1201 = s_1164[1:0];
  assign s_1202 = s_1128[1:0];
  assign s_1203 = s_1204[3];
  assign s_1204 = {s_1205,s_1275};
  assign s_1205 = s_1206 & s_1241;
  assign s_1206 = s_1207[2];
  assign s_1207 = {s_1208,s_1235};
  assign s_1208 = s_1209 & s_1223;
  assign s_1209 = s_1210[1];
  assign s_1210 = {s_1211,s_1219};
  assign s_1211 = s_1212 & s_1217;
  assign s_1212 = ~s_1213;
  assign s_1213 = s_1214[1];
  assign s_1214 = s_1215[3:2];
  assign s_1215 = s_1216[7:4];
  assign s_1216 = s_1138[7:0];
  assign s_1217 = ~s_1218;
  assign s_1218 = s_1214[0];
  assign s_1219 = s_1220 & s_1222;
  assign s_1220 = ~s_1221;
  assign s_1221 = s_1214[1];
  assign s_1222 = s_1214[0];
  assign s_1223 = s_1224[1];
  assign s_1224 = {s_1225,s_1231};
  assign s_1225 = s_1226 & s_1229;
  assign s_1226 = ~s_1227;
  assign s_1227 = s_1228[1];
  assign s_1228 = s_1215[1:0];
  assign s_1229 = ~s_1230;
  assign s_1230 = s_1228[0];
  assign s_1231 = s_1232 & s_1234;
  assign s_1232 = ~s_1233;
  assign s_1233 = s_1228[1];
  assign s_1234 = s_1228[0];
  assign s_1235 = {s_1236,s_1238};
  assign s_1236 = s_1209 & s_1237;
  assign s_1237 = ~s_1223;
  assign s_1238 = s_1209?s_1239:s_1240;
  assign s_1239 = s_1224[0:0];
  assign s_1240 = s_1210[0:0];
  assign s_1241 = s_1242[2];
  assign s_1242 = {s_1243,s_1269};
  assign s_1243 = s_1244 & s_1257;
  assign s_1244 = s_1245[1];
  assign s_1245 = {s_1246,s_1253};
  assign s_1246 = s_1247 & s_1251;
  assign s_1247 = ~s_1248;
  assign s_1248 = s_1249[1];
  assign s_1249 = s_1250[3:2];
  assign s_1250 = s_1216[3:0];
  assign s_1251 = ~s_1252;
  assign s_1252 = s_1249[0];
  assign s_1253 = s_1254 & s_1256;
  assign s_1254 = ~s_1255;
  assign s_1255 = s_1249[1];
  assign s_1256 = s_1249[0];
  assign s_1257 = s_1258[1];
  assign s_1258 = {s_1259,s_1265};
  assign s_1259 = s_1260 & s_1263;
  assign s_1260 = ~s_1261;
  assign s_1261 = s_1262[1];
  assign s_1262 = s_1250[1:0];
  assign s_1263 = ~s_1264;
  assign s_1264 = s_1262[0];
  assign s_1265 = s_1266 & s_1268;
  assign s_1266 = ~s_1267;
  assign s_1267 = s_1262[1];
  assign s_1268 = s_1262[0];
  assign s_1269 = {s_1270,s_1272};
  assign s_1270 = s_1244 & s_1271;
  assign s_1271 = ~s_1257;
  assign s_1272 = s_1244?s_1273:s_1274;
  assign s_1273 = s_1258[0:0];
  assign s_1274 = s_1245[0:0];
  assign s_1275 = {s_1276,s_1278};
  assign s_1276 = s_1206 & s_1277;
  assign s_1277 = ~s_1241;
  assign s_1278 = s_1206?s_1279:s_1280;
  assign s_1279 = s_1242[1:0];
  assign s_1280 = s_1207[1:0];
  assign s_1281 = {s_1282,s_1284};
  assign s_1282 = s_1124 & s_1283;
  assign s_1283 = ~s_1203;
  assign s_1284 = s_1124?s_1285:s_1286;
  assign s_1285 = s_1204[2:0];
  assign s_1286 = s_1125[2:0];
  assign s_1287 = {s_1288,s_1290};
  assign s_1288 = s_953 & s_1289;
  assign s_1289 = ~s_1121;
  assign s_1290 = s_953?s_1291:s_1292;
  assign s_1291 = s_1122[3:0];
  assign s_1292 = s_954[3:0];
  assign s_1293 = s_1294[5];
  assign s_1294 = {s_1295,s_1629};
  assign s_1295 = s_1296 & s_1463;
  assign s_1296 = s_1297[4];
  assign s_1297 = {s_1298,s_1457};
  assign s_1298 = s_1299 & s_1379;
  assign s_1299 = s_1300[3];
  assign s_1300 = {s_1301,s_1373};
  assign s_1301 = s_1302 & s_1339;
  assign s_1302 = s_1303[2];
  assign s_1303 = {s_1304,s_1333};
  assign s_1304 = s_1305 & s_1321;
  assign s_1305 = s_1306[1];
  assign s_1306 = {s_1307,s_1317};
  assign s_1307 = s_1308 & s_1315;
  assign s_1308 = ~s_1309;
  assign s_1309 = s_1310[1];
  assign s_1310 = s_1311[3:2];
  assign s_1311 = s_1312[7:4];
  assign s_1312 = s_1313[15:8];
  assign s_1313 = s_1314[31:16];
  assign s_1314 = s_972[31:0];
  assign s_1315 = ~s_1316;
  assign s_1316 = s_1310[0];
  assign s_1317 = s_1318 & s_1320;
  assign s_1318 = ~s_1319;
  assign s_1319 = s_1310[1];
  assign s_1320 = s_1310[0];
  assign s_1321 = s_1322[1];
  assign s_1322 = {s_1323,s_1329};
  assign s_1323 = s_1324 & s_1327;
  assign s_1324 = ~s_1325;
  assign s_1325 = s_1326[1];
  assign s_1326 = s_1311[1:0];
  assign s_1327 = ~s_1328;
  assign s_1328 = s_1326[0];
  assign s_1329 = s_1330 & s_1332;
  assign s_1330 = ~s_1331;
  assign s_1331 = s_1326[1];
  assign s_1332 = s_1326[0];
  assign s_1333 = {s_1334,s_1336};
  assign s_1334 = s_1305 & s_1335;
  assign s_1335 = ~s_1321;
  assign s_1336 = s_1305?s_1337:s_1338;
  assign s_1337 = s_1322[0:0];
  assign s_1338 = s_1306[0:0];
  assign s_1339 = s_1340[2];
  assign s_1340 = {s_1341,s_1367};
  assign s_1341 = s_1342 & s_1355;
  assign s_1342 = s_1343[1];
  assign s_1343 = {s_1344,s_1351};
  assign s_1344 = s_1345 & s_1349;
  assign s_1345 = ~s_1346;
  assign s_1346 = s_1347[1];
  assign s_1347 = s_1348[3:2];
  assign s_1348 = s_1312[3:0];
  assign s_1349 = ~s_1350;
  assign s_1350 = s_1347[0];
  assign s_1351 = s_1352 & s_1354;
  assign s_1352 = ~s_1353;
  assign s_1353 = s_1347[1];
  assign s_1354 = s_1347[0];
  assign s_1355 = s_1356[1];
  assign s_1356 = {s_1357,s_1363};
  assign s_1357 = s_1358 & s_1361;
  assign s_1358 = ~s_1359;
  assign s_1359 = s_1360[1];
  assign s_1360 = s_1348[1:0];
  assign s_1361 = ~s_1362;
  assign s_1362 = s_1360[0];
  assign s_1363 = s_1364 & s_1366;
  assign s_1364 = ~s_1365;
  assign s_1365 = s_1360[1];
  assign s_1366 = s_1360[0];
  assign s_1367 = {s_1368,s_1370};
  assign s_1368 = s_1342 & s_1369;
  assign s_1369 = ~s_1355;
  assign s_1370 = s_1342?s_1371:s_1372;
  assign s_1371 = s_1356[0:0];
  assign s_1372 = s_1343[0:0];
  assign s_1373 = {s_1374,s_1376};
  assign s_1374 = s_1302 & s_1375;
  assign s_1375 = ~s_1339;
  assign s_1376 = s_1302?s_1377:s_1378;
  assign s_1377 = s_1340[1:0];
  assign s_1378 = s_1303[1:0];
  assign s_1379 = s_1380[3];
  assign s_1380 = {s_1381,s_1451};
  assign s_1381 = s_1382 & s_1417;
  assign s_1382 = s_1383[2];
  assign s_1383 = {s_1384,s_1411};
  assign s_1384 = s_1385 & s_1399;
  assign s_1385 = s_1386[1];
  assign s_1386 = {s_1387,s_1395};
  assign s_1387 = s_1388 & s_1393;
  assign s_1388 = ~s_1389;
  assign s_1389 = s_1390[1];
  assign s_1390 = s_1391[3:2];
  assign s_1391 = s_1392[7:4];
  assign s_1392 = s_1313[7:0];
  assign s_1393 = ~s_1394;
  assign s_1394 = s_1390[0];
  assign s_1395 = s_1396 & s_1398;
  assign s_1396 = ~s_1397;
  assign s_1397 = s_1390[1];
  assign s_1398 = s_1390[0];
  assign s_1399 = s_1400[1];
  assign s_1400 = {s_1401,s_1407};
  assign s_1401 = s_1402 & s_1405;
  assign s_1402 = ~s_1403;
  assign s_1403 = s_1404[1];
  assign s_1404 = s_1391[1:0];
  assign s_1405 = ~s_1406;
  assign s_1406 = s_1404[0];
  assign s_1407 = s_1408 & s_1410;
  assign s_1408 = ~s_1409;
  assign s_1409 = s_1404[1];
  assign s_1410 = s_1404[0];
  assign s_1411 = {s_1412,s_1414};
  assign s_1412 = s_1385 & s_1413;
  assign s_1413 = ~s_1399;
  assign s_1414 = s_1385?s_1415:s_1416;
  assign s_1415 = s_1400[0:0];
  assign s_1416 = s_1386[0:0];
  assign s_1417 = s_1418[2];
  assign s_1418 = {s_1419,s_1445};
  assign s_1419 = s_1420 & s_1433;
  assign s_1420 = s_1421[1];
  assign s_1421 = {s_1422,s_1429};
  assign s_1422 = s_1423 & s_1427;
  assign s_1423 = ~s_1424;
  assign s_1424 = s_1425[1];
  assign s_1425 = s_1426[3:2];
  assign s_1426 = s_1392[3:0];
  assign s_1427 = ~s_1428;
  assign s_1428 = s_1425[0];
  assign s_1429 = s_1430 & s_1432;
  assign s_1430 = ~s_1431;
  assign s_1431 = s_1425[1];
  assign s_1432 = s_1425[0];
  assign s_1433 = s_1434[1];
  assign s_1434 = {s_1435,s_1441};
  assign s_1435 = s_1436 & s_1439;
  assign s_1436 = ~s_1437;
  assign s_1437 = s_1438[1];
  assign s_1438 = s_1426[1:0];
  assign s_1439 = ~s_1440;
  assign s_1440 = s_1438[0];
  assign s_1441 = s_1442 & s_1444;
  assign s_1442 = ~s_1443;
  assign s_1443 = s_1438[1];
  assign s_1444 = s_1438[0];
  assign s_1445 = {s_1446,s_1448};
  assign s_1446 = s_1420 & s_1447;
  assign s_1447 = ~s_1433;
  assign s_1448 = s_1420?s_1449:s_1450;
  assign s_1449 = s_1434[0:0];
  assign s_1450 = s_1421[0:0];
  assign s_1451 = {s_1452,s_1454};
  assign s_1452 = s_1382 & s_1453;
  assign s_1453 = ~s_1417;
  assign s_1454 = s_1382?s_1455:s_1456;
  assign s_1455 = s_1418[1:0];
  assign s_1456 = s_1383[1:0];
  assign s_1457 = {s_1458,s_1460};
  assign s_1458 = s_1299 & s_1459;
  assign s_1459 = ~s_1379;
  assign s_1460 = s_1299?s_1461:s_1462;
  assign s_1461 = s_1380[2:0];
  assign s_1462 = s_1300[2:0];
  assign s_1463 = s_1464[4];
  assign s_1464 = {s_1465,s_1623};
  assign s_1465 = s_1466 & s_1545;
  assign s_1466 = s_1467[3];
  assign s_1467 = {s_1468,s_1539};
  assign s_1468 = s_1469 & s_1505;
  assign s_1469 = s_1470[2];
  assign s_1470 = {s_1471,s_1499};
  assign s_1471 = s_1472 & s_1487;
  assign s_1472 = s_1473[1];
  assign s_1473 = {s_1474,s_1483};
  assign s_1474 = s_1475 & s_1481;
  assign s_1475 = ~s_1476;
  assign s_1476 = s_1477[1];
  assign s_1477 = s_1478[3:2];
  assign s_1478 = s_1479[7:4];
  assign s_1479 = s_1480[15:8];
  assign s_1480 = s_1314[15:0];
  assign s_1481 = ~s_1482;
  assign s_1482 = s_1477[0];
  assign s_1483 = s_1484 & s_1486;
  assign s_1484 = ~s_1485;
  assign s_1485 = s_1477[1];
  assign s_1486 = s_1477[0];
  assign s_1487 = s_1488[1];
  assign s_1488 = {s_1489,s_1495};
  assign s_1489 = s_1490 & s_1493;
  assign s_1490 = ~s_1491;
  assign s_1491 = s_1492[1];
  assign s_1492 = s_1478[1:0];
  assign s_1493 = ~s_1494;
  assign s_1494 = s_1492[0];
  assign s_1495 = s_1496 & s_1498;
  assign s_1496 = ~s_1497;
  assign s_1497 = s_1492[1];
  assign s_1498 = s_1492[0];
  assign s_1499 = {s_1500,s_1502};
  assign s_1500 = s_1472 & s_1501;
  assign s_1501 = ~s_1487;
  assign s_1502 = s_1472?s_1503:s_1504;
  assign s_1503 = s_1488[0:0];
  assign s_1504 = s_1473[0:0];
  assign s_1505 = s_1506[2];
  assign s_1506 = {s_1507,s_1533};
  assign s_1507 = s_1508 & s_1521;
  assign s_1508 = s_1509[1];
  assign s_1509 = {s_1510,s_1517};
  assign s_1510 = s_1511 & s_1515;
  assign s_1511 = ~s_1512;
  assign s_1512 = s_1513[1];
  assign s_1513 = s_1514[3:2];
  assign s_1514 = s_1479[3:0];
  assign s_1515 = ~s_1516;
  assign s_1516 = s_1513[0];
  assign s_1517 = s_1518 & s_1520;
  assign s_1518 = ~s_1519;
  assign s_1519 = s_1513[1];
  assign s_1520 = s_1513[0];
  assign s_1521 = s_1522[1];
  assign s_1522 = {s_1523,s_1529};
  assign s_1523 = s_1524 & s_1527;
  assign s_1524 = ~s_1525;
  assign s_1525 = s_1526[1];
  assign s_1526 = s_1514[1:0];
  assign s_1527 = ~s_1528;
  assign s_1528 = s_1526[0];
  assign s_1529 = s_1530 & s_1532;
  assign s_1530 = ~s_1531;
  assign s_1531 = s_1526[1];
  assign s_1532 = s_1526[0];
  assign s_1533 = {s_1534,s_1536};
  assign s_1534 = s_1508 & s_1535;
  assign s_1535 = ~s_1521;
  assign s_1536 = s_1508?s_1537:s_1538;
  assign s_1537 = s_1522[0:0];
  assign s_1538 = s_1509[0:0];
  assign s_1539 = {s_1540,s_1542};
  assign s_1540 = s_1469 & s_1541;
  assign s_1541 = ~s_1505;
  assign s_1542 = s_1469?s_1543:s_1544;
  assign s_1543 = s_1506[1:0];
  assign s_1544 = s_1470[1:0];
  assign s_1545 = s_1546[3];
  assign s_1546 = {s_1547,s_1617};
  assign s_1547 = s_1548 & s_1583;
  assign s_1548 = s_1549[2];
  assign s_1549 = {s_1550,s_1577};
  assign s_1550 = s_1551 & s_1565;
  assign s_1551 = s_1552[1];
  assign s_1552 = {s_1553,s_1561};
  assign s_1553 = s_1554 & s_1559;
  assign s_1554 = ~s_1555;
  assign s_1555 = s_1556[1];
  assign s_1556 = s_1557[3:2];
  assign s_1557 = s_1558[7:4];
  assign s_1558 = s_1480[7:0];
  assign s_1559 = ~s_1560;
  assign s_1560 = s_1556[0];
  assign s_1561 = s_1562 & s_1564;
  assign s_1562 = ~s_1563;
  assign s_1563 = s_1556[1];
  assign s_1564 = s_1556[0];
  assign s_1565 = s_1566[1];
  assign s_1566 = {s_1567,s_1573};
  assign s_1567 = s_1568 & s_1571;
  assign s_1568 = ~s_1569;
  assign s_1569 = s_1570[1];
  assign s_1570 = s_1557[1:0];
  assign s_1571 = ~s_1572;
  assign s_1572 = s_1570[0];
  assign s_1573 = s_1574 & s_1576;
  assign s_1574 = ~s_1575;
  assign s_1575 = s_1570[1];
  assign s_1576 = s_1570[0];
  assign s_1577 = {s_1578,s_1580};
  assign s_1578 = s_1551 & s_1579;
  assign s_1579 = ~s_1565;
  assign s_1580 = s_1551?s_1581:s_1582;
  assign s_1581 = s_1566[0:0];
  assign s_1582 = s_1552[0:0];
  assign s_1583 = s_1584[2];
  assign s_1584 = {s_1585,s_1611};
  assign s_1585 = s_1586 & s_1599;
  assign s_1586 = s_1587[1];
  assign s_1587 = {s_1588,s_1595};
  assign s_1588 = s_1589 & s_1593;
  assign s_1589 = ~s_1590;
  assign s_1590 = s_1591[1];
  assign s_1591 = s_1592[3:2];
  assign s_1592 = s_1558[3:0];
  assign s_1593 = ~s_1594;
  assign s_1594 = s_1591[0];
  assign s_1595 = s_1596 & s_1598;
  assign s_1596 = ~s_1597;
  assign s_1597 = s_1591[1];
  assign s_1598 = s_1591[0];
  assign s_1599 = s_1600[1];
  assign s_1600 = {s_1601,s_1607};
  assign s_1601 = s_1602 & s_1605;
  assign s_1602 = ~s_1603;
  assign s_1603 = s_1604[1];
  assign s_1604 = s_1592[1:0];
  assign s_1605 = ~s_1606;
  assign s_1606 = s_1604[0];
  assign s_1607 = s_1608 & s_1610;
  assign s_1608 = ~s_1609;
  assign s_1609 = s_1604[1];
  assign s_1610 = s_1604[0];
  assign s_1611 = {s_1612,s_1614};
  assign s_1612 = s_1586 & s_1613;
  assign s_1613 = ~s_1599;
  assign s_1614 = s_1586?s_1615:s_1616;
  assign s_1615 = s_1600[0:0];
  assign s_1616 = s_1587[0:0];
  assign s_1617 = {s_1618,s_1620};
  assign s_1618 = s_1548 & s_1619;
  assign s_1619 = ~s_1583;
  assign s_1620 = s_1548?s_1621:s_1622;
  assign s_1621 = s_1584[1:0];
  assign s_1622 = s_1549[1:0];
  assign s_1623 = {s_1624,s_1626};
  assign s_1624 = s_1466 & s_1625;
  assign s_1625 = ~s_1545;
  assign s_1626 = s_1466?s_1627:s_1628;
  assign s_1627 = s_1546[2:0];
  assign s_1628 = s_1467[2:0];
  assign s_1629 = {s_1630,s_1632};
  assign s_1630 = s_1296 & s_1631;
  assign s_1631 = ~s_1463;
  assign s_1632 = s_1296?s_1633:s_1634;
  assign s_1633 = s_1464[3:0];
  assign s_1634 = s_1297[3:0];
  assign s_1635 = {s_1636,s_1638};
  assign s_1636 = s_950 & s_1637;
  assign s_1637 = ~s_1293;
  assign s_1638 = s_950?s_1639:s_1640;
  assign s_1639 = s_1294[4:0];
  assign s_1640 = s_951[4:0];
  assign s_1641 = {s_1642,s_1644};
  assign s_1642 = s_209 & s_1643;
  assign s_1643 = ~s_947;
  assign s_1644 = s_209?s_1645:s_1646;
  assign s_1645 = s_948[5:0];
  assign s_1646 = s_210[5:0];
  dq #(13, 16) dq_s_1647 (clk, s_1647, s_1648);
  assign s_1648 = s_1649 - s_1651;
  dq #(13, 1) dq_s_1649 (clk, s_1649, s_1650);
  assign s_1650 = s_194 + s_190;
  assign s_1651 = -13'd1022;
  assign s_1652 = s_1653 <= s_1654;
  assign s_1653 = s_206;
  dq #(13, 16) dq_s_1654 (clk, s_1654, s_1648);
  assign s_1655 = 1'd1;
  dq #(53, 1) dq_s_1656 (clk, s_1656, s_30);
  assign s_1657 = s_1658 & s_1660;
  dq #(1, 1) dq_s_1658 (clk, s_1658, s_1659);
  assign s_1659 = s_31[52];
  assign s_1660 = s_1661 | s_1668;
  assign s_1661 = s_1662 | s_1664;
  dq #(1, 1) dq_s_1662 (clk, s_1662, s_1663);
  assign s_1663 = s_31[51];
  dq #(1, 1) dq_s_1664 (clk, s_1664, s_1665);
  assign s_1665 = s_1666 != s_1667;
  assign s_1666 = s_31[50:0];
  assign s_1667 = 53'd0;
  dq #(1, 1) dq_s_1668 (clk, s_1668, s_1669);
  assign s_1669 = s_30[0];
  assign s_1670 = s_26[52:0];
  assign s_1671 = s_26[53];
  assign s_1672 = {s_1673,s_1684};
  assign s_1673 = {s_1674,s_1675};
  dq #(1, 21) dq_s_1674 (clk, s_1674, s_3);
  assign s_1675 = s_1676 + s_1683;
  assign s_1676 = s_1677[10:0];
  dq #(13, 1) dq_s_1677 (clk, s_1677, s_1678);
  assign s_1678 = s_1679 + s_1671;
  dq #(13, 1) dq_s_1679 (clk, s_1679, s_1680);
  dq #(13, 1) dq_s_1680 (clk, s_1680, s_1681);
  assign s_1681 = s_1682 - s_204;
  dq #(13, 17) dq_s_1682 (clk, s_1682, s_1649);
  assign s_1683 = 10'd1023;
  assign s_1684 = s_23[51:0];
  assign s_1685 = s_1686 & s_1688;
  assign s_1686 = s_1676 == s_1687;
  assign s_1687 = -11'd1022;
  assign s_1688 = ~s_1689;
  assign s_1689 = s_23[52];
  assign s_1690 = s_23 == s_1691;
  assign s_1691 = 53'd0;
  assign s_1692 = s_1693 | s_1702;
  assign s_1693 = s_1694 | s_1696;
  assign s_1694 = $signed(s_1677) > $signed(s_1695);
  assign s_1695 = 12'd1023;
  dq #(1, 21) dq_s_1696 (clk, s_1696, s_1697);
  assign s_1697 = s_1698 & s_1700;
  assign s_1698 = s_52 == s_1699;
  assign s_1699 = 11'd1024;
  assign s_1700 = s_56 == s_1701;
  assign s_1701 = 52'd0;
  dq #(1, 21) dq_s_1702 (clk, s_1702, s_1703);
  assign s_1703 = s_1704 & s_1706;
  assign s_1704 = s_64 == s_1705;
  assign s_1705 = 11'd1024;
  assign s_1706 = s_68 == s_1707;
  assign s_1707 = 52'd0;
  dq #(1, 21) dq_s_1708 (clk, s_1708, s_1709);
  assign s_1709 = s_1710 | s_1715;
  assign s_1710 = s_1711 & s_1713;
  assign s_1711 = s_52 == s_1712;
  assign s_1712 = 11'd1024;
  assign s_1713 = s_56 != s_1714;
  assign s_1714 = 52'd0;
  assign s_1715 = s_1716 & s_1718;
  assign s_1716 = s_64 == s_1717;
  assign s_1717 = 11'd1024;
  assign s_1718 = s_68 != s_1719;
  assign s_1719 = 52'd0;
  assign double_mul_z = s_0;
endmodule
