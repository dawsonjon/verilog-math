module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module sqrt(clk, sqrt_a, sqrt_z);
  input clk;
  input [31:0] sqrt_a;
  output [31:0] sqrt_z;
  wire [31:0] s_0;
  wire [31:0] s_1;
  wire [31:0] s_2;
  wire [0:0] s_3;
  wire [31:0] s_4;
  wire [30:0] s_5;
  wire [31:0] s_6;
  wire [31:0] s_7;
  wire [31:0] s_8;
  wire [30:0] s_9;
  wire [31:0] s_10;
  wire [31:0] s_11;
  wire [31:0] s_12;
  wire [30:0] s_13;
  wire [31:0] s_14;
  wire [31:0] s_15;
  wire [8:0] s_16;
  wire [8:0] s_17;
  wire [7:0] s_18;
  wire [22:0] s_19;
  wire [23:0] s_20;
  wire [23:0] s_21;
  wire [23:0] s_22;
  wire [24:0] s_23;
  wire [24:0] s_24;
  wire [24:0] s_25;
  wire [23:0] s_26;
  wire [24:0] s_27;
  wire [24:0] s_28;
  wire [24:0] s_29;
  wire [24:0] s_30;
  wire [24:0] s_31;
  wire [24:0] s_32;
  wire [24:0] s_33;
  wire [50:0] s_34;
  wire [50:0] s_35;
  wire [50:0] s_36;
  wire [50:0] s_37;
  wire [50:0] s_38;
  wire [50:0] s_39;
  wire [50:0] s_40;
  wire [50:0] s_41;
  wire [50:0] s_42;
  wire [50:0] s_43;
  wire [50:0] s_44;
  wire [50:0] s_45;
  wire [50:0] s_46;
  wire [50:0] s_47;
  wire [50:0] s_48;
  wire [50:0] s_49;
  wire [50:0] s_50;
  wire [50:0] s_51;
  wire [50:0] s_52;
  wire [50:0] s_53;
  wire [50:0] s_54;
  wire [50:0] s_55;
  wire [50:0] s_56;
  wire [50:0] s_57;
  wire [50:0] s_58;
  wire [50:0] s_59;
  wire [50:0] s_60;
  wire [50:0] s_61;
  wire [50:0] s_62;
  wire [50:0] s_63;
  wire [50:0] s_64;
  wire [50:0] s_65;
  wire [50:0] s_66;
  wire [50:0] s_67;
  wire [50:0] s_68;
  wire [50:0] s_69;
  wire [50:0] s_70;
  wire [50:0] s_71;
  wire [50:0] s_72;
  wire [50:0] s_73;
  wire [50:0] s_74;
  wire [50:0] s_75;
  wire [50:0] s_76;
  wire [50:0] s_77;
  wire [50:0] s_78;
  wire [50:0] s_79;
  wire [50:0] s_80;
  wire [50:0] s_81;
  wire [50:0] s_82;
  wire [50:0] s_83;
  wire [50:0] s_84;
  wire [50:0] s_85;
  wire [50:0] s_86;
  wire [25:0] s_87;
  wire [50:0] s_88;
  wire [0:0] s_89;
  wire [51:0] s_90;
  wire [51:0] s_91;
  wire [51:0] s_92;
  wire [51:0] s_93;
  wire [25:0] s_94;
  wire [4:0] s_95;
  wire [50:0] s_96;
  wire [50:0] s_97;
  wire [50:0] s_98;
  wire [50:0] s_99;
  wire [50:0] s_100;
  wire [23:0] s_101;
  wire [23:0] s_102;
  wire [23:0] s_103;
  wire [23:0] s_104;
  wire [0:0] s_105;
  wire [0:0] s_106;
  wire [0:0] s_107;
  wire [0:0] s_108;
  wire [7:0] s_109;
  wire [7:0] s_110;
  wire [6:0] s_111;
  wire [7:0] s_112;
  wire [22:0] s_113;
  wire [9:0] s_114;
  wire [9:0] s_115;
  wire [5:0] s_116;
  wire [5:0] s_117;
  wire [0:0] s_118;
  wire [0:0] s_119;
  wire [4:0] s_120;
  wire [0:0] s_121;
  wire [0:0] s_122;
  wire [3:0] s_123;
  wire [0:0] s_124;
  wire [0:0] s_125;
  wire [2:0] s_126;
  wire [0:0] s_127;
  wire [0:0] s_128;
  wire [1:0] s_129;
  wire [0:0] s_130;
  wire [0:0] s_131;
  wire [0:0] s_132;
  wire [1:0] s_133;
  wire [3:0] s_134;
  wire [7:0] s_135;
  wire [15:0] s_136;
  wire [31:0] s_137;
  wire [30:0] s_138;
  wire [29:0] s_139;
  wire [28:0] s_140;
  wire [27:0] s_141;
  wire [26:0] s_142;
  wire [25:0] s_143;
  wire [24:0] s_144;
  wire [0:0] s_145;
  wire [0:0] s_146;
  wire [0:0] s_147;
  wire [0:0] s_148;
  wire [0:0] s_149;
  wire [0:0] s_150;
  wire [0:0] s_151;
  wire [0:0] s_152;
  wire [0:0] s_153;
  wire [0:0] s_154;
  wire [0:0] s_155;
  wire [0:0] s_156;
  wire [0:0] s_157;
  wire [0:0] s_158;
  wire [0:0] s_159;
  wire [1:0] s_160;
  wire [0:0] s_161;
  wire [0:0] s_162;
  wire [0:0] s_163;
  wire [1:0] s_164;
  wire [0:0] s_165;
  wire [0:0] s_166;
  wire [0:0] s_167;
  wire [0:0] s_168;
  wire [0:0] s_169;
  wire [0:0] s_170;
  wire [1:0] s_171;
  wire [0:0] s_172;
  wire [0:0] s_173;
  wire [0:0] s_174;
  wire [0:0] s_175;
  wire [0:0] s_176;
  wire [0:0] s_177;
  wire [2:0] s_178;
  wire [0:0] s_179;
  wire [0:0] s_180;
  wire [1:0] s_181;
  wire [0:0] s_182;
  wire [0:0] s_183;
  wire [0:0] s_184;
  wire [1:0] s_185;
  wire [3:0] s_186;
  wire [0:0] s_187;
  wire [0:0] s_188;
  wire [0:0] s_189;
  wire [0:0] s_190;
  wire [0:0] s_191;
  wire [0:0] s_192;
  wire [0:0] s_193;
  wire [1:0] s_194;
  wire [0:0] s_195;
  wire [0:0] s_196;
  wire [0:0] s_197;
  wire [1:0] s_198;
  wire [0:0] s_199;
  wire [0:0] s_200;
  wire [0:0] s_201;
  wire [0:0] s_202;
  wire [0:0] s_203;
  wire [0:0] s_204;
  wire [1:0] s_205;
  wire [0:0] s_206;
  wire [0:0] s_207;
  wire [0:0] s_208;
  wire [0:0] s_209;
  wire [0:0] s_210;
  wire [2:0] s_211;
  wire [0:0] s_212;
  wire [0:0] s_213;
  wire [1:0] s_214;
  wire [1:0] s_215;
  wire [1:0] s_216;
  wire [0:0] s_217;
  wire [3:0] s_218;
  wire [0:0] s_219;
  wire [0:0] s_220;
  wire [2:0] s_221;
  wire [0:0] s_222;
  wire [0:0] s_223;
  wire [1:0] s_224;
  wire [0:0] s_225;
  wire [0:0] s_226;
  wire [0:0] s_227;
  wire [1:0] s_228;
  wire [3:0] s_229;
  wire [7:0] s_230;
  wire [0:0] s_231;
  wire [0:0] s_232;
  wire [0:0] s_233;
  wire [0:0] s_234;
  wire [0:0] s_235;
  wire [0:0] s_236;
  wire [0:0] s_237;
  wire [1:0] s_238;
  wire [0:0] s_239;
  wire [0:0] s_240;
  wire [0:0] s_241;
  wire [1:0] s_242;
  wire [0:0] s_243;
  wire [0:0] s_244;
  wire [0:0] s_245;
  wire [0:0] s_246;
  wire [0:0] s_247;
  wire [0:0] s_248;
  wire [1:0] s_249;
  wire [0:0] s_250;
  wire [0:0] s_251;
  wire [0:0] s_252;
  wire [0:0] s_253;
  wire [0:0] s_254;
  wire [0:0] s_255;
  wire [2:0] s_256;
  wire [0:0] s_257;
  wire [0:0] s_258;
  wire [1:0] s_259;
  wire [0:0] s_260;
  wire [0:0] s_261;
  wire [0:0] s_262;
  wire [1:0] s_263;
  wire [3:0] s_264;
  wire [0:0] s_265;
  wire [0:0] s_266;
  wire [0:0] s_267;
  wire [0:0] s_268;
  wire [0:0] s_269;
  wire [0:0] s_270;
  wire [0:0] s_271;
  wire [1:0] s_272;
  wire [0:0] s_273;
  wire [0:0] s_274;
  wire [0:0] s_275;
  wire [1:0] s_276;
  wire [0:0] s_277;
  wire [0:0] s_278;
  wire [0:0] s_279;
  wire [0:0] s_280;
  wire [0:0] s_281;
  wire [0:0] s_282;
  wire [1:0] s_283;
  wire [0:0] s_284;
  wire [0:0] s_285;
  wire [0:0] s_286;
  wire [0:0] s_287;
  wire [0:0] s_288;
  wire [2:0] s_289;
  wire [0:0] s_290;
  wire [0:0] s_291;
  wire [1:0] s_292;
  wire [1:0] s_293;
  wire [1:0] s_294;
  wire [3:0] s_295;
  wire [0:0] s_296;
  wire [0:0] s_297;
  wire [2:0] s_298;
  wire [2:0] s_299;
  wire [2:0] s_300;
  wire [0:0] s_301;
  wire [4:0] s_302;
  wire [0:0] s_303;
  wire [0:0] s_304;
  wire [3:0] s_305;
  wire [0:0] s_306;
  wire [0:0] s_307;
  wire [2:0] s_308;
  wire [0:0] s_309;
  wire [0:0] s_310;
  wire [1:0] s_311;
  wire [0:0] s_312;
  wire [0:0] s_313;
  wire [0:0] s_314;
  wire [1:0] s_315;
  wire [3:0] s_316;
  wire [7:0] s_317;
  wire [15:0] s_318;
  wire [0:0] s_319;
  wire [0:0] s_320;
  wire [0:0] s_321;
  wire [0:0] s_322;
  wire [0:0] s_323;
  wire [0:0] s_324;
  wire [0:0] s_325;
  wire [1:0] s_326;
  wire [0:0] s_327;
  wire [0:0] s_328;
  wire [0:0] s_329;
  wire [1:0] s_330;
  wire [0:0] s_331;
  wire [0:0] s_332;
  wire [0:0] s_333;
  wire [0:0] s_334;
  wire [0:0] s_335;
  wire [0:0] s_336;
  wire [1:0] s_337;
  wire [0:0] s_338;
  wire [0:0] s_339;
  wire [0:0] s_340;
  wire [0:0] s_341;
  wire [0:0] s_342;
  wire [0:0] s_343;
  wire [2:0] s_344;
  wire [0:0] s_345;
  wire [0:0] s_346;
  wire [1:0] s_347;
  wire [0:0] s_348;
  wire [0:0] s_349;
  wire [0:0] s_350;
  wire [1:0] s_351;
  wire [3:0] s_352;
  wire [0:0] s_353;
  wire [0:0] s_354;
  wire [0:0] s_355;
  wire [0:0] s_356;
  wire [0:0] s_357;
  wire [0:0] s_358;
  wire [0:0] s_359;
  wire [1:0] s_360;
  wire [0:0] s_361;
  wire [0:0] s_362;
  wire [0:0] s_363;
  wire [1:0] s_364;
  wire [0:0] s_365;
  wire [0:0] s_366;
  wire [0:0] s_367;
  wire [0:0] s_368;
  wire [0:0] s_369;
  wire [0:0] s_370;
  wire [1:0] s_371;
  wire [0:0] s_372;
  wire [0:0] s_373;
  wire [0:0] s_374;
  wire [0:0] s_375;
  wire [0:0] s_376;
  wire [2:0] s_377;
  wire [0:0] s_378;
  wire [0:0] s_379;
  wire [1:0] s_380;
  wire [1:0] s_381;
  wire [1:0] s_382;
  wire [0:0] s_383;
  wire [3:0] s_384;
  wire [0:0] s_385;
  wire [0:0] s_386;
  wire [2:0] s_387;
  wire [0:0] s_388;
  wire [0:0] s_389;
  wire [1:0] s_390;
  wire [0:0] s_391;
  wire [0:0] s_392;
  wire [0:0] s_393;
  wire [1:0] s_394;
  wire [3:0] s_395;
  wire [7:0] s_396;
  wire [0:0] s_397;
  wire [0:0] s_398;
  wire [0:0] s_399;
  wire [0:0] s_400;
  wire [0:0] s_401;
  wire [0:0] s_402;
  wire [0:0] s_403;
  wire [1:0] s_404;
  wire [0:0] s_405;
  wire [0:0] s_406;
  wire [0:0] s_407;
  wire [1:0] s_408;
  wire [0:0] s_409;
  wire [0:0] s_410;
  wire [0:0] s_411;
  wire [0:0] s_412;
  wire [0:0] s_413;
  wire [0:0] s_414;
  wire [1:0] s_415;
  wire [0:0] s_416;
  wire [0:0] s_417;
  wire [0:0] s_418;
  wire [0:0] s_419;
  wire [0:0] s_420;
  wire [0:0] s_421;
  wire [2:0] s_422;
  wire [0:0] s_423;
  wire [0:0] s_424;
  wire [1:0] s_425;
  wire [0:0] s_426;
  wire [0:0] s_427;
  wire [0:0] s_428;
  wire [1:0] s_429;
  wire [3:0] s_430;
  wire [0:0] s_431;
  wire [0:0] s_432;
  wire [0:0] s_433;
  wire [0:0] s_434;
  wire [0:0] s_435;
  wire [0:0] s_436;
  wire [0:0] s_437;
  wire [1:0] s_438;
  wire [0:0] s_439;
  wire [0:0] s_440;
  wire [0:0] s_441;
  wire [1:0] s_442;
  wire [0:0] s_443;
  wire [0:0] s_444;
  wire [0:0] s_445;
  wire [0:0] s_446;
  wire [0:0] s_447;
  wire [0:0] s_448;
  wire [1:0] s_449;
  wire [0:0] s_450;
  wire [0:0] s_451;
  wire [0:0] s_452;
  wire [0:0] s_453;
  wire [0:0] s_454;
  wire [2:0] s_455;
  wire [0:0] s_456;
  wire [0:0] s_457;
  wire [1:0] s_458;
  wire [1:0] s_459;
  wire [1:0] s_460;
  wire [3:0] s_461;
  wire [0:0] s_462;
  wire [0:0] s_463;
  wire [2:0] s_464;
  wire [2:0] s_465;
  wire [2:0] s_466;
  wire [4:0] s_467;
  wire [0:0] s_468;
  wire [0:0] s_469;
  wire [3:0] s_470;
  wire [3:0] s_471;
  wire [3:0] s_472;
  wire [9:0] s_473;
  wire [9:0] s_474;
  wire [9:0] s_475;
  wire [7:0] s_476;
  wire [7:0] s_477;
  wire [9:0] s_478;
  wire [0:0] s_479;
  wire [9:0] s_480;
  wire [9:0] s_481;
  wire [0:0] s_482;
  wire [0:0] s_483;
  wire [9:0] s_484;
  wire [9:0] s_485;
  wire [9:0] s_486;
  wire [4:0] s_487;
  wire [50:0] s_488;
  wire [0:0] s_489;
  wire [51:0] s_490;
  wire [51:0] s_491;
  wire [51:0] s_492;
  wire [51:0] s_493;
  wire [50:0] s_494;
  wire [4:0] s_495;
  wire [48:0] s_496;
  wire [50:0] s_497;
  wire [0:0] s_498;
  wire [51:0] s_499;
  wire [51:0] s_500;
  wire [51:0] s_501;
  wire [50:0] s_502;
  wire [4:0] s_503;
  wire [46:0] s_504;
  wire [50:0] s_505;
  wire [0:0] s_506;
  wire [51:0] s_507;
  wire [51:0] s_508;
  wire [51:0] s_509;
  wire [50:0] s_510;
  wire [4:0] s_511;
  wire [44:0] s_512;
  wire [50:0] s_513;
  wire [0:0] s_514;
  wire [51:0] s_515;
  wire [51:0] s_516;
  wire [51:0] s_517;
  wire [50:0] s_518;
  wire [4:0] s_519;
  wire [42:0] s_520;
  wire [50:0] s_521;
  wire [0:0] s_522;
  wire [51:0] s_523;
  wire [51:0] s_524;
  wire [51:0] s_525;
  wire [50:0] s_526;
  wire [4:0] s_527;
  wire [40:0] s_528;
  wire [50:0] s_529;
  wire [0:0] s_530;
  wire [51:0] s_531;
  wire [51:0] s_532;
  wire [51:0] s_533;
  wire [50:0] s_534;
  wire [4:0] s_535;
  wire [38:0] s_536;
  wire [50:0] s_537;
  wire [0:0] s_538;
  wire [51:0] s_539;
  wire [51:0] s_540;
  wire [51:0] s_541;
  wire [50:0] s_542;
  wire [4:0] s_543;
  wire [36:0] s_544;
  wire [50:0] s_545;
  wire [0:0] s_546;
  wire [51:0] s_547;
  wire [51:0] s_548;
  wire [51:0] s_549;
  wire [50:0] s_550;
  wire [4:0] s_551;
  wire [34:0] s_552;
  wire [50:0] s_553;
  wire [0:0] s_554;
  wire [51:0] s_555;
  wire [51:0] s_556;
  wire [51:0] s_557;
  wire [50:0] s_558;
  wire [4:0] s_559;
  wire [32:0] s_560;
  wire [50:0] s_561;
  wire [0:0] s_562;
  wire [51:0] s_563;
  wire [51:0] s_564;
  wire [51:0] s_565;
  wire [50:0] s_566;
  wire [4:0] s_567;
  wire [30:0] s_568;
  wire [50:0] s_569;
  wire [0:0] s_570;
  wire [51:0] s_571;
  wire [51:0] s_572;
  wire [51:0] s_573;
  wire [50:0] s_574;
  wire [3:0] s_575;
  wire [28:0] s_576;
  wire [50:0] s_577;
  wire [0:0] s_578;
  wire [51:0] s_579;
  wire [51:0] s_580;
  wire [51:0] s_581;
  wire [50:0] s_582;
  wire [3:0] s_583;
  wire [26:0] s_584;
  wire [50:0] s_585;
  wire [0:0] s_586;
  wire [51:0] s_587;
  wire [51:0] s_588;
  wire [51:0] s_589;
  wire [50:0] s_590;
  wire [3:0] s_591;
  wire [24:0] s_592;
  wire [50:0] s_593;
  wire [0:0] s_594;
  wire [51:0] s_595;
  wire [51:0] s_596;
  wire [51:0] s_597;
  wire [50:0] s_598;
  wire [3:0] s_599;
  wire [22:0] s_600;
  wire [50:0] s_601;
  wire [0:0] s_602;
  wire [51:0] s_603;
  wire [51:0] s_604;
  wire [51:0] s_605;
  wire [50:0] s_606;
  wire [3:0] s_607;
  wire [20:0] s_608;
  wire [50:0] s_609;
  wire [0:0] s_610;
  wire [51:0] s_611;
  wire [51:0] s_612;
  wire [51:0] s_613;
  wire [50:0] s_614;
  wire [3:0] s_615;
  wire [18:0] s_616;
  wire [50:0] s_617;
  wire [0:0] s_618;
  wire [51:0] s_619;
  wire [51:0] s_620;
  wire [51:0] s_621;
  wire [50:0] s_622;
  wire [3:0] s_623;
  wire [16:0] s_624;
  wire [50:0] s_625;
  wire [0:0] s_626;
  wire [51:0] s_627;
  wire [51:0] s_628;
  wire [51:0] s_629;
  wire [50:0] s_630;
  wire [3:0] s_631;
  wire [14:0] s_632;
  wire [50:0] s_633;
  wire [0:0] s_634;
  wire [51:0] s_635;
  wire [51:0] s_636;
  wire [51:0] s_637;
  wire [50:0] s_638;
  wire [2:0] s_639;
  wire [12:0] s_640;
  wire [50:0] s_641;
  wire [0:0] s_642;
  wire [51:0] s_643;
  wire [51:0] s_644;
  wire [51:0] s_645;
  wire [50:0] s_646;
  wire [2:0] s_647;
  wire [10:0] s_648;
  wire [50:0] s_649;
  wire [0:0] s_650;
  wire [51:0] s_651;
  wire [51:0] s_652;
  wire [51:0] s_653;
  wire [50:0] s_654;
  wire [2:0] s_655;
  wire [8:0] s_656;
  wire [50:0] s_657;
  wire [0:0] s_658;
  wire [51:0] s_659;
  wire [51:0] s_660;
  wire [51:0] s_661;
  wire [50:0] s_662;
  wire [2:0] s_663;
  wire [6:0] s_664;
  wire [50:0] s_665;
  wire [0:0] s_666;
  wire [51:0] s_667;
  wire [51:0] s_668;
  wire [51:0] s_669;
  wire [50:0] s_670;
  wire [1:0] s_671;
  wire [4:0] s_672;
  wire [50:0] s_673;
  wire [0:0] s_674;
  wire [51:0] s_675;
  wire [51:0] s_676;
  wire [51:0] s_677;
  wire [50:0] s_678;
  wire [1:0] s_679;
  wire [2:0] s_680;
  wire [50:0] s_681;
  wire [0:0] s_682;
  wire [51:0] s_683;
  wire [51:0] s_684;
  wire [51:0] s_685;
  wire [50:0] s_686;
  wire [0:0] s_687;
  wire [0:0] s_688;
  wire [9:0] s_689;
  wire [9:0] s_690;
  wire [0:0] s_691;
  wire [9:0] s_692;
  wire [9:0] s_693;
  wire [9:0] s_694;
  wire [9:0] s_695;
  wire [9:0] s_696;
  wire [9:0] s_697;
  wire [0:0] s_698;
  wire [9:0] s_699;
  wire [0:0] s_700;
  wire [9:0] s_701;
  wire [9:0] s_702;
  wire [5:0] s_703;
  wire [5:0] s_704;
  wire [0:0] s_705;
  wire [0:0] s_706;
  wire [4:0] s_707;
  wire [0:0] s_708;
  wire [0:0] s_709;
  wire [3:0] s_710;
  wire [0:0] s_711;
  wire [0:0] s_712;
  wire [2:0] s_713;
  wire [0:0] s_714;
  wire [0:0] s_715;
  wire [1:0] s_716;
  wire [0:0] s_717;
  wire [0:0] s_718;
  wire [0:0] s_719;
  wire [1:0] s_720;
  wire [3:0] s_721;
  wire [7:0] s_722;
  wire [15:0] s_723;
  wire [31:0] s_724;
  wire [30:0] s_725;
  wire [29:0] s_726;
  wire [28:0] s_727;
  wire [27:0] s_728;
  wire [26:0] s_729;
  wire [25:0] s_730;
  wire [0:0] s_731;
  wire [0:0] s_732;
  wire [0:0] s_733;
  wire [0:0] s_734;
  wire [0:0] s_735;
  wire [0:0] s_736;
  wire [0:0] s_737;
  wire [0:0] s_738;
  wire [0:0] s_739;
  wire [0:0] s_740;
  wire [0:0] s_741;
  wire [0:0] s_742;
  wire [0:0] s_743;
  wire [0:0] s_744;
  wire [1:0] s_745;
  wire [0:0] s_746;
  wire [0:0] s_747;
  wire [0:0] s_748;
  wire [1:0] s_749;
  wire [0:0] s_750;
  wire [0:0] s_751;
  wire [0:0] s_752;
  wire [0:0] s_753;
  wire [0:0] s_754;
  wire [0:0] s_755;
  wire [1:0] s_756;
  wire [0:0] s_757;
  wire [0:0] s_758;
  wire [0:0] s_759;
  wire [0:0] s_760;
  wire [0:0] s_761;
  wire [0:0] s_762;
  wire [2:0] s_763;
  wire [0:0] s_764;
  wire [0:0] s_765;
  wire [1:0] s_766;
  wire [0:0] s_767;
  wire [0:0] s_768;
  wire [0:0] s_769;
  wire [1:0] s_770;
  wire [3:0] s_771;
  wire [0:0] s_772;
  wire [0:0] s_773;
  wire [0:0] s_774;
  wire [0:0] s_775;
  wire [0:0] s_776;
  wire [0:0] s_777;
  wire [0:0] s_778;
  wire [1:0] s_779;
  wire [0:0] s_780;
  wire [0:0] s_781;
  wire [0:0] s_782;
  wire [1:0] s_783;
  wire [0:0] s_784;
  wire [0:0] s_785;
  wire [0:0] s_786;
  wire [0:0] s_787;
  wire [0:0] s_788;
  wire [0:0] s_789;
  wire [1:0] s_790;
  wire [0:0] s_791;
  wire [0:0] s_792;
  wire [0:0] s_793;
  wire [0:0] s_794;
  wire [0:0] s_795;
  wire [2:0] s_796;
  wire [0:0] s_797;
  wire [0:0] s_798;
  wire [1:0] s_799;
  wire [1:0] s_800;
  wire [1:0] s_801;
  wire [0:0] s_802;
  wire [3:0] s_803;
  wire [0:0] s_804;
  wire [0:0] s_805;
  wire [2:0] s_806;
  wire [0:0] s_807;
  wire [0:0] s_808;
  wire [1:0] s_809;
  wire [0:0] s_810;
  wire [0:0] s_811;
  wire [0:0] s_812;
  wire [1:0] s_813;
  wire [3:0] s_814;
  wire [7:0] s_815;
  wire [0:0] s_816;
  wire [0:0] s_817;
  wire [0:0] s_818;
  wire [0:0] s_819;
  wire [0:0] s_820;
  wire [0:0] s_821;
  wire [0:0] s_822;
  wire [1:0] s_823;
  wire [0:0] s_824;
  wire [0:0] s_825;
  wire [0:0] s_826;
  wire [1:0] s_827;
  wire [0:0] s_828;
  wire [0:0] s_829;
  wire [0:0] s_830;
  wire [0:0] s_831;
  wire [0:0] s_832;
  wire [0:0] s_833;
  wire [1:0] s_834;
  wire [0:0] s_835;
  wire [0:0] s_836;
  wire [0:0] s_837;
  wire [0:0] s_838;
  wire [0:0] s_839;
  wire [0:0] s_840;
  wire [2:0] s_841;
  wire [0:0] s_842;
  wire [0:0] s_843;
  wire [1:0] s_844;
  wire [0:0] s_845;
  wire [0:0] s_846;
  wire [0:0] s_847;
  wire [1:0] s_848;
  wire [3:0] s_849;
  wire [0:0] s_850;
  wire [0:0] s_851;
  wire [0:0] s_852;
  wire [0:0] s_853;
  wire [0:0] s_854;
  wire [0:0] s_855;
  wire [0:0] s_856;
  wire [1:0] s_857;
  wire [0:0] s_858;
  wire [0:0] s_859;
  wire [0:0] s_860;
  wire [1:0] s_861;
  wire [0:0] s_862;
  wire [0:0] s_863;
  wire [0:0] s_864;
  wire [0:0] s_865;
  wire [0:0] s_866;
  wire [0:0] s_867;
  wire [1:0] s_868;
  wire [0:0] s_869;
  wire [0:0] s_870;
  wire [0:0] s_871;
  wire [0:0] s_872;
  wire [0:0] s_873;
  wire [2:0] s_874;
  wire [0:0] s_875;
  wire [0:0] s_876;
  wire [1:0] s_877;
  wire [1:0] s_878;
  wire [1:0] s_879;
  wire [3:0] s_880;
  wire [0:0] s_881;
  wire [0:0] s_882;
  wire [2:0] s_883;
  wire [2:0] s_884;
  wire [2:0] s_885;
  wire [0:0] s_886;
  wire [4:0] s_887;
  wire [0:0] s_888;
  wire [0:0] s_889;
  wire [3:0] s_890;
  wire [0:0] s_891;
  wire [0:0] s_892;
  wire [2:0] s_893;
  wire [0:0] s_894;
  wire [0:0] s_895;
  wire [1:0] s_896;
  wire [0:0] s_897;
  wire [0:0] s_898;
  wire [0:0] s_899;
  wire [1:0] s_900;
  wire [3:0] s_901;
  wire [7:0] s_902;
  wire [15:0] s_903;
  wire [0:0] s_904;
  wire [0:0] s_905;
  wire [0:0] s_906;
  wire [0:0] s_907;
  wire [0:0] s_908;
  wire [0:0] s_909;
  wire [0:0] s_910;
  wire [1:0] s_911;
  wire [0:0] s_912;
  wire [0:0] s_913;
  wire [0:0] s_914;
  wire [1:0] s_915;
  wire [0:0] s_916;
  wire [0:0] s_917;
  wire [0:0] s_918;
  wire [0:0] s_919;
  wire [0:0] s_920;
  wire [0:0] s_921;
  wire [1:0] s_922;
  wire [0:0] s_923;
  wire [0:0] s_924;
  wire [0:0] s_925;
  wire [0:0] s_926;
  wire [0:0] s_927;
  wire [0:0] s_928;
  wire [2:0] s_929;
  wire [0:0] s_930;
  wire [0:0] s_931;
  wire [1:0] s_932;
  wire [0:0] s_933;
  wire [0:0] s_934;
  wire [0:0] s_935;
  wire [1:0] s_936;
  wire [3:0] s_937;
  wire [0:0] s_938;
  wire [0:0] s_939;
  wire [0:0] s_940;
  wire [0:0] s_941;
  wire [0:0] s_942;
  wire [0:0] s_943;
  wire [0:0] s_944;
  wire [1:0] s_945;
  wire [0:0] s_946;
  wire [0:0] s_947;
  wire [0:0] s_948;
  wire [1:0] s_949;
  wire [0:0] s_950;
  wire [0:0] s_951;
  wire [0:0] s_952;
  wire [0:0] s_953;
  wire [0:0] s_954;
  wire [0:0] s_955;
  wire [1:0] s_956;
  wire [0:0] s_957;
  wire [0:0] s_958;
  wire [0:0] s_959;
  wire [0:0] s_960;
  wire [0:0] s_961;
  wire [2:0] s_962;
  wire [0:0] s_963;
  wire [0:0] s_964;
  wire [1:0] s_965;
  wire [1:0] s_966;
  wire [1:0] s_967;
  wire [0:0] s_968;
  wire [3:0] s_969;
  wire [0:0] s_970;
  wire [0:0] s_971;
  wire [2:0] s_972;
  wire [0:0] s_973;
  wire [0:0] s_974;
  wire [1:0] s_975;
  wire [0:0] s_976;
  wire [0:0] s_977;
  wire [0:0] s_978;
  wire [1:0] s_979;
  wire [3:0] s_980;
  wire [7:0] s_981;
  wire [0:0] s_982;
  wire [0:0] s_983;
  wire [0:0] s_984;
  wire [0:0] s_985;
  wire [0:0] s_986;
  wire [0:0] s_987;
  wire [0:0] s_988;
  wire [1:0] s_989;
  wire [0:0] s_990;
  wire [0:0] s_991;
  wire [0:0] s_992;
  wire [1:0] s_993;
  wire [0:0] s_994;
  wire [0:0] s_995;
  wire [0:0] s_996;
  wire [0:0] s_997;
  wire [0:0] s_998;
  wire [0:0] s_999;
  wire [1:0] s_1000;
  wire [0:0] s_1001;
  wire [0:0] s_1002;
  wire [0:0] s_1003;
  wire [0:0] s_1004;
  wire [0:0] s_1005;
  wire [0:0] s_1006;
  wire [2:0] s_1007;
  wire [0:0] s_1008;
  wire [0:0] s_1009;
  wire [1:0] s_1010;
  wire [0:0] s_1011;
  wire [0:0] s_1012;
  wire [0:0] s_1013;
  wire [1:0] s_1014;
  wire [3:0] s_1015;
  wire [0:0] s_1016;
  wire [0:0] s_1017;
  wire [0:0] s_1018;
  wire [0:0] s_1019;
  wire [0:0] s_1020;
  wire [0:0] s_1021;
  wire [0:0] s_1022;
  wire [1:0] s_1023;
  wire [0:0] s_1024;
  wire [0:0] s_1025;
  wire [0:0] s_1026;
  wire [1:0] s_1027;
  wire [0:0] s_1028;
  wire [0:0] s_1029;
  wire [0:0] s_1030;
  wire [0:0] s_1031;
  wire [0:0] s_1032;
  wire [0:0] s_1033;
  wire [1:0] s_1034;
  wire [0:0] s_1035;
  wire [0:0] s_1036;
  wire [0:0] s_1037;
  wire [0:0] s_1038;
  wire [0:0] s_1039;
  wire [2:0] s_1040;
  wire [0:0] s_1041;
  wire [0:0] s_1042;
  wire [1:0] s_1043;
  wire [1:0] s_1044;
  wire [1:0] s_1045;
  wire [3:0] s_1046;
  wire [0:0] s_1047;
  wire [0:0] s_1048;
  wire [2:0] s_1049;
  wire [2:0] s_1050;
  wire [2:0] s_1051;
  wire [4:0] s_1052;
  wire [0:0] s_1053;
  wire [0:0] s_1054;
  wire [3:0] s_1055;
  wire [3:0] s_1056;
  wire [3:0] s_1057;
  wire [9:0] s_1058;
  wire [9:0] s_1059;
  wire [9:0] s_1060;
  wire [9:0] s_1061;
  wire [9:0] s_1062;
  wire [9:0] s_1063;
  wire [0:0] s_1064;
  wire [9:0] s_1065;
  wire [9:0] s_1066;
  wire [0:0] s_1067;
  wire [0:0] s_1068;
  wire [0:0] s_1069;
  wire [0:0] s_1070;
  wire [0:0] s_1071;
  wire [0:0] s_1072;
  wire [0:0] s_1073;
  wire [0:0] s_1074;
  wire [0:0] s_1075;
  wire [23:0] s_1076;
  wire [0:0] s_1077;
  wire [31:0] s_1078;
  wire [8:0] s_1079;
  wire [0:0] s_1080;
  wire [7:0] s_1081;
  wire [7:0] s_1082;
  wire [9:0] s_1083;
  wire [9:0] s_1084;
  wire [9:0] s_1085;
  wire [9:0] s_1086;
  wire [9:0] s_1087;
  wire [6:0] s_1088;
  wire [22:0] s_1089;
  wire [0:0] s_1090;
  wire [0:0] s_1091;
  wire [7:0] s_1092;
  wire [0:0] s_1093;
  wire [0:0] s_1094;
  wire [0:0] s_1095;
  wire [23:0] s_1096;
  wire [0:0] s_1097;
  wire [0:0] s_1098;
  wire [0:0] s_1099;
  wire [7:0] s_1100;
  wire [0:0] s_1101;
  wire [22:0] s_1102;
  wire [0:0] s_1103;
  wire [0:0] s_1104;
  wire [0:0] s_1105;
  wire [0:0] s_1106;
  wire [7:0] s_1107;
  wire [0:0] s_1108;
  wire [22:0] s_1109;
  wire [0:0] s_1110;
  wire [0:0] s_1111;
  wire [0:0] s_1112;
  wire [0:0] s_1113;

  assign s_0 = s_1103?s_1:s_6;
  dq #(32, 10) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_5};
  assign s_3 = s_4[31];
  assign s_4 = sqrt_a;
  assign s_5 = 31'd2143289344;
  assign s_6 = s_1097?s_7:s_10;
  dq #(32, 10) dq_s_7 (clk, s_7, s_8);
  assign s_8 = {s_3,s_9};
  assign s_9 = 31'd2139095040;
  assign s_10 = s_1095?s_11:s_14;
  dq #(32, 10) dq_s_11 (clk, s_11, s_12);
  assign s_12 = {s_3,s_13};
  assign s_13 = 31'd0;
  assign s_14 = s_1090?s_15:s_1078;
  assign s_15 = {s_16,s_19};
  dq #(9, 10) dq_s_16 (clk, s_16, s_17);
  assign s_17 = {s_3,s_18};
  assign s_18 = 8'd0;
  assign s_19 = s_20[22:0];
  dq #(24, 1) dq_s_20 (clk, s_20, s_21);
  assign s_21 = s_1077?s_22:s_1076;
  assign s_22 = s_23[24:1];
  assign s_23 = s_1068?s_24:s_26;
  assign s_24 = s_25 + s_1067;
  assign s_25 = s_26;
  assign s_26 = s_27[24:1];
  dq #(25, 1) dq_s_27 (clk, s_27, s_28);
  assign s_28 = s_29 << s_701;
  dq #(25, 2) dq_s_29 (clk, s_29, s_30);
  dq #(25, 1) dq_s_30 (clk, s_30, s_31);
  assign s_31 = s_32 >> s_689;
  dq #(25, 2) dq_s_32 (clk, s_32, s_33);
  assign s_33 = s_34[24:0];
  assign s_34 = s_682?s_35:s_36;
  assign s_35 = s_36 + s_681;
  assign s_36 = s_674?s_37:s_38;
  assign s_37 = s_38 + s_673;
  assign s_38 = s_666?s_39:s_40;
  assign s_39 = s_40 + s_665;
  assign s_40 = s_658?s_41:s_42;
  assign s_41 = s_42 + s_657;
  assign s_42 = s_650?s_43:s_44;
  assign s_43 = s_44 + s_649;
  assign s_44 = s_642?s_45:s_46;
  assign s_45 = s_46 + s_641;
  assign s_46 = s_634?s_47:s_48;
  assign s_47 = s_48 + s_633;
  assign s_48 = s_626?s_49:s_50;
  assign s_49 = s_50 + s_625;
  assign s_50 = s_618?s_51:s_52;
  assign s_51 = s_52 + s_617;
  assign s_52 = s_610?s_53:s_54;
  assign s_53 = s_54 + s_609;
  assign s_54 = s_602?s_55:s_56;
  assign s_55 = s_56 + s_601;
  assign s_56 = s_594?s_57:s_58;
  assign s_57 = s_58 + s_593;
  assign s_58 = s_586?s_59:s_60;
  assign s_59 = s_60 + s_585;
  assign s_60 = s_578?s_61:s_62;
  assign s_61 = s_62 + s_577;
  assign s_62 = s_570?s_63:s_64;
  assign s_63 = s_64 + s_569;
  assign s_64 = s_562?s_65:s_66;
  assign s_65 = s_66 + s_561;
  assign s_66 = s_554?s_67:s_68;
  assign s_67 = s_68 + s_553;
  assign s_68 = s_546?s_69:s_70;
  assign s_69 = s_70 + s_545;
  assign s_70 = s_538?s_71:s_72;
  assign s_71 = s_72 + s_537;
  assign s_72 = s_530?s_73:s_74;
  assign s_73 = s_74 + s_529;
  assign s_74 = s_522?s_75:s_76;
  assign s_75 = s_76 + s_521;
  assign s_76 = s_514?s_77:s_78;
  assign s_77 = s_78 + s_513;
  assign s_78 = s_506?s_79:s_80;
  assign s_79 = s_80 + s_505;
  assign s_80 = s_498?s_81:s_82;
  assign s_81 = s_82 + s_497;
  assign s_82 = s_489?s_83:s_84;
  assign s_83 = s_84 + s_488;
  assign s_84 = s_89?s_85:s_87;
  dq #(51, 3) dq_s_85 (clk, s_85, s_86);
  assign s_86 = s_87 + s_88;
  assign s_87 = 26'd0;
  assign s_88 = 51'd33554432;
  assign s_89 = s_90 <= s_97;
  dq #(52, 3) dq_s_90 (clk, s_90, s_91);
  assign s_91 = s_92 | s_96;
  assign s_92 = s_93 + s_94;
  assign s_93 = 52'd0;
  assign s_94 = s_87 << s_95;
  assign s_95 = 5'd26;
  assign s_96 = 51'd1125899906842624;
  assign s_97 = s_98 << s_487;
  assign s_98 = s_483?s_99:s_100;
  assign s_99 = s_100 << s_482;
  assign s_100 = s_101;
  dq #(24, 1) dq_s_101 (clk, s_101, s_102);
  assign s_102 = s_103 << s_114;
  dq #(24, 2) dq_s_103 (clk, s_103, s_104);
  assign s_104 = {s_105,s_113};
  assign s_105 = s_108?s_106:s_107;
  assign s_106 = 1'd0;
  assign s_107 = 1'd1;
  assign s_108 = s_109 == s_112;
  assign s_109 = s_110 - s_111;
  assign s_110 = s_4[30:23];
  assign s_111 = 7'd127;
  assign s_112 = -8'd127;
  assign s_113 = s_4[22:0];
  dq #(10, 1) dq_s_114 (clk, s_114, s_115);
  assign s_115 = s_479?s_116:s_473;
  dq #(6, 1) dq_s_116 (clk, s_116, s_117);
  assign s_117 = {s_118,s_467};
  assign s_118 = s_119 & s_301;
  assign s_119 = s_120[4];
  assign s_120 = {s_121,s_295};
  assign s_121 = s_122 & s_217;
  assign s_122 = s_123[3];
  assign s_123 = {s_124,s_211};
  assign s_124 = s_125 & s_177;
  assign s_125 = s_126[2];
  assign s_126 = {s_127,s_171};
  assign s_127 = s_128 & s_159;
  assign s_128 = s_129[1];
  assign s_129 = {s_130,s_155};
  assign s_130 = s_131 & s_153;
  assign s_131 = ~s_132;
  assign s_132 = s_133[1];
  assign s_133 = s_134[3:2];
  assign s_134 = s_135[7:4];
  assign s_135 = s_136[15:8];
  assign s_136 = s_137[31:16];
  assign s_137 = {s_138,s_152};
  assign s_138 = {s_139,s_151};
  assign s_139 = {s_140,s_150};
  assign s_140 = {s_141,s_149};
  assign s_141 = {s_142,s_148};
  assign s_142 = {s_143,s_147};
  assign s_143 = {s_144,s_146};
  assign s_144 = {s_104,s_145};
  assign s_145 = 1'd1;
  assign s_146 = 1'd1;
  assign s_147 = 1'd1;
  assign s_148 = 1'd1;
  assign s_149 = 1'd1;
  assign s_150 = 1'd1;
  assign s_151 = 1'd1;
  assign s_152 = 1'd1;
  assign s_153 = ~s_154;
  assign s_154 = s_133[0];
  assign s_155 = s_156 & s_158;
  assign s_156 = ~s_157;
  assign s_157 = s_133[1];
  assign s_158 = s_133[0];
  assign s_159 = s_160[1];
  assign s_160 = {s_161,s_167};
  assign s_161 = s_162 & s_165;
  assign s_162 = ~s_163;
  assign s_163 = s_164[1];
  assign s_164 = s_134[1:0];
  assign s_165 = ~s_166;
  assign s_166 = s_164[0];
  assign s_167 = s_168 & s_170;
  assign s_168 = ~s_169;
  assign s_169 = s_164[1];
  assign s_170 = s_164[0];
  assign s_171 = {s_172,s_174};
  assign s_172 = s_128 & s_173;
  assign s_173 = ~s_159;
  assign s_174 = s_128?s_175:s_176;
  assign s_175 = s_160[0:0];
  assign s_176 = s_129[0:0];
  assign s_177 = s_178[2];
  assign s_178 = {s_179,s_205};
  assign s_179 = s_180 & s_193;
  assign s_180 = s_181[1];
  assign s_181 = {s_182,s_189};
  assign s_182 = s_183 & s_187;
  assign s_183 = ~s_184;
  assign s_184 = s_185[1];
  assign s_185 = s_186[3:2];
  assign s_186 = s_135[3:0];
  assign s_187 = ~s_188;
  assign s_188 = s_185[0];
  assign s_189 = s_190 & s_192;
  assign s_190 = ~s_191;
  assign s_191 = s_185[1];
  assign s_192 = s_185[0];
  assign s_193 = s_194[1];
  assign s_194 = {s_195,s_201};
  assign s_195 = s_196 & s_199;
  assign s_196 = ~s_197;
  assign s_197 = s_198[1];
  assign s_198 = s_186[1:0];
  assign s_199 = ~s_200;
  assign s_200 = s_198[0];
  assign s_201 = s_202 & s_204;
  assign s_202 = ~s_203;
  assign s_203 = s_198[1];
  assign s_204 = s_198[0];
  assign s_205 = {s_206,s_208};
  assign s_206 = s_180 & s_207;
  assign s_207 = ~s_193;
  assign s_208 = s_180?s_209:s_210;
  assign s_209 = s_194[0:0];
  assign s_210 = s_181[0:0];
  assign s_211 = {s_212,s_214};
  assign s_212 = s_125 & s_213;
  assign s_213 = ~s_177;
  assign s_214 = s_125?s_215:s_216;
  assign s_215 = s_178[1:0];
  assign s_216 = s_126[1:0];
  assign s_217 = s_218[3];
  assign s_218 = {s_219,s_289};
  assign s_219 = s_220 & s_255;
  assign s_220 = s_221[2];
  assign s_221 = {s_222,s_249};
  assign s_222 = s_223 & s_237;
  assign s_223 = s_224[1];
  assign s_224 = {s_225,s_233};
  assign s_225 = s_226 & s_231;
  assign s_226 = ~s_227;
  assign s_227 = s_228[1];
  assign s_228 = s_229[3:2];
  assign s_229 = s_230[7:4];
  assign s_230 = s_136[7:0];
  assign s_231 = ~s_232;
  assign s_232 = s_228[0];
  assign s_233 = s_234 & s_236;
  assign s_234 = ~s_235;
  assign s_235 = s_228[1];
  assign s_236 = s_228[0];
  assign s_237 = s_238[1];
  assign s_238 = {s_239,s_245};
  assign s_239 = s_240 & s_243;
  assign s_240 = ~s_241;
  assign s_241 = s_242[1];
  assign s_242 = s_229[1:0];
  assign s_243 = ~s_244;
  assign s_244 = s_242[0];
  assign s_245 = s_246 & s_248;
  assign s_246 = ~s_247;
  assign s_247 = s_242[1];
  assign s_248 = s_242[0];
  assign s_249 = {s_250,s_252};
  assign s_250 = s_223 & s_251;
  assign s_251 = ~s_237;
  assign s_252 = s_223?s_253:s_254;
  assign s_253 = s_238[0:0];
  assign s_254 = s_224[0:0];
  assign s_255 = s_256[2];
  assign s_256 = {s_257,s_283};
  assign s_257 = s_258 & s_271;
  assign s_258 = s_259[1];
  assign s_259 = {s_260,s_267};
  assign s_260 = s_261 & s_265;
  assign s_261 = ~s_262;
  assign s_262 = s_263[1];
  assign s_263 = s_264[3:2];
  assign s_264 = s_230[3:0];
  assign s_265 = ~s_266;
  assign s_266 = s_263[0];
  assign s_267 = s_268 & s_270;
  assign s_268 = ~s_269;
  assign s_269 = s_263[1];
  assign s_270 = s_263[0];
  assign s_271 = s_272[1];
  assign s_272 = {s_273,s_279};
  assign s_273 = s_274 & s_277;
  assign s_274 = ~s_275;
  assign s_275 = s_276[1];
  assign s_276 = s_264[1:0];
  assign s_277 = ~s_278;
  assign s_278 = s_276[0];
  assign s_279 = s_280 & s_282;
  assign s_280 = ~s_281;
  assign s_281 = s_276[1];
  assign s_282 = s_276[0];
  assign s_283 = {s_284,s_286};
  assign s_284 = s_258 & s_285;
  assign s_285 = ~s_271;
  assign s_286 = s_258?s_287:s_288;
  assign s_287 = s_272[0:0];
  assign s_288 = s_259[0:0];
  assign s_289 = {s_290,s_292};
  assign s_290 = s_220 & s_291;
  assign s_291 = ~s_255;
  assign s_292 = s_220?s_293:s_294;
  assign s_293 = s_256[1:0];
  assign s_294 = s_221[1:0];
  assign s_295 = {s_296,s_298};
  assign s_296 = s_122 & s_297;
  assign s_297 = ~s_217;
  assign s_298 = s_122?s_299:s_300;
  assign s_299 = s_218[2:0];
  assign s_300 = s_123[2:0];
  assign s_301 = s_302[4];
  assign s_302 = {s_303,s_461};
  assign s_303 = s_304 & s_383;
  assign s_304 = s_305[3];
  assign s_305 = {s_306,s_377};
  assign s_306 = s_307 & s_343;
  assign s_307 = s_308[2];
  assign s_308 = {s_309,s_337};
  assign s_309 = s_310 & s_325;
  assign s_310 = s_311[1];
  assign s_311 = {s_312,s_321};
  assign s_312 = s_313 & s_319;
  assign s_313 = ~s_314;
  assign s_314 = s_315[1];
  assign s_315 = s_316[3:2];
  assign s_316 = s_317[7:4];
  assign s_317 = s_318[15:8];
  assign s_318 = s_137[15:0];
  assign s_319 = ~s_320;
  assign s_320 = s_315[0];
  assign s_321 = s_322 & s_324;
  assign s_322 = ~s_323;
  assign s_323 = s_315[1];
  assign s_324 = s_315[0];
  assign s_325 = s_326[1];
  assign s_326 = {s_327,s_333};
  assign s_327 = s_328 & s_331;
  assign s_328 = ~s_329;
  assign s_329 = s_330[1];
  assign s_330 = s_316[1:0];
  assign s_331 = ~s_332;
  assign s_332 = s_330[0];
  assign s_333 = s_334 & s_336;
  assign s_334 = ~s_335;
  assign s_335 = s_330[1];
  assign s_336 = s_330[0];
  assign s_337 = {s_338,s_340};
  assign s_338 = s_310 & s_339;
  assign s_339 = ~s_325;
  assign s_340 = s_310?s_341:s_342;
  assign s_341 = s_326[0:0];
  assign s_342 = s_311[0:0];
  assign s_343 = s_344[2];
  assign s_344 = {s_345,s_371};
  assign s_345 = s_346 & s_359;
  assign s_346 = s_347[1];
  assign s_347 = {s_348,s_355};
  assign s_348 = s_349 & s_353;
  assign s_349 = ~s_350;
  assign s_350 = s_351[1];
  assign s_351 = s_352[3:2];
  assign s_352 = s_317[3:0];
  assign s_353 = ~s_354;
  assign s_354 = s_351[0];
  assign s_355 = s_356 & s_358;
  assign s_356 = ~s_357;
  assign s_357 = s_351[1];
  assign s_358 = s_351[0];
  assign s_359 = s_360[1];
  assign s_360 = {s_361,s_367};
  assign s_361 = s_362 & s_365;
  assign s_362 = ~s_363;
  assign s_363 = s_364[1];
  assign s_364 = s_352[1:0];
  assign s_365 = ~s_366;
  assign s_366 = s_364[0];
  assign s_367 = s_368 & s_370;
  assign s_368 = ~s_369;
  assign s_369 = s_364[1];
  assign s_370 = s_364[0];
  assign s_371 = {s_372,s_374};
  assign s_372 = s_346 & s_373;
  assign s_373 = ~s_359;
  assign s_374 = s_346?s_375:s_376;
  assign s_375 = s_360[0:0];
  assign s_376 = s_347[0:0];
  assign s_377 = {s_378,s_380};
  assign s_378 = s_307 & s_379;
  assign s_379 = ~s_343;
  assign s_380 = s_307?s_381:s_382;
  assign s_381 = s_344[1:0];
  assign s_382 = s_308[1:0];
  assign s_383 = s_384[3];
  assign s_384 = {s_385,s_455};
  assign s_385 = s_386 & s_421;
  assign s_386 = s_387[2];
  assign s_387 = {s_388,s_415};
  assign s_388 = s_389 & s_403;
  assign s_389 = s_390[1];
  assign s_390 = {s_391,s_399};
  assign s_391 = s_392 & s_397;
  assign s_392 = ~s_393;
  assign s_393 = s_394[1];
  assign s_394 = s_395[3:2];
  assign s_395 = s_396[7:4];
  assign s_396 = s_318[7:0];
  assign s_397 = ~s_398;
  assign s_398 = s_394[0];
  assign s_399 = s_400 & s_402;
  assign s_400 = ~s_401;
  assign s_401 = s_394[1];
  assign s_402 = s_394[0];
  assign s_403 = s_404[1];
  assign s_404 = {s_405,s_411};
  assign s_405 = s_406 & s_409;
  assign s_406 = ~s_407;
  assign s_407 = s_408[1];
  assign s_408 = s_395[1:0];
  assign s_409 = ~s_410;
  assign s_410 = s_408[0];
  assign s_411 = s_412 & s_414;
  assign s_412 = ~s_413;
  assign s_413 = s_408[1];
  assign s_414 = s_408[0];
  assign s_415 = {s_416,s_418};
  assign s_416 = s_389 & s_417;
  assign s_417 = ~s_403;
  assign s_418 = s_389?s_419:s_420;
  assign s_419 = s_404[0:0];
  assign s_420 = s_390[0:0];
  assign s_421 = s_422[2];
  assign s_422 = {s_423,s_449};
  assign s_423 = s_424 & s_437;
  assign s_424 = s_425[1];
  assign s_425 = {s_426,s_433};
  assign s_426 = s_427 & s_431;
  assign s_427 = ~s_428;
  assign s_428 = s_429[1];
  assign s_429 = s_430[3:2];
  assign s_430 = s_396[3:0];
  assign s_431 = ~s_432;
  assign s_432 = s_429[0];
  assign s_433 = s_434 & s_436;
  assign s_434 = ~s_435;
  assign s_435 = s_429[1];
  assign s_436 = s_429[0];
  assign s_437 = s_438[1];
  assign s_438 = {s_439,s_445};
  assign s_439 = s_440 & s_443;
  assign s_440 = ~s_441;
  assign s_441 = s_442[1];
  assign s_442 = s_430[1:0];
  assign s_443 = ~s_444;
  assign s_444 = s_442[0];
  assign s_445 = s_446 & s_448;
  assign s_446 = ~s_447;
  assign s_447 = s_442[1];
  assign s_448 = s_442[0];
  assign s_449 = {s_450,s_452};
  assign s_450 = s_424 & s_451;
  assign s_451 = ~s_437;
  assign s_452 = s_424?s_453:s_454;
  assign s_453 = s_438[0:0];
  assign s_454 = s_425[0:0];
  assign s_455 = {s_456,s_458};
  assign s_456 = s_386 & s_457;
  assign s_457 = ~s_421;
  assign s_458 = s_386?s_459:s_460;
  assign s_459 = s_422[1:0];
  assign s_460 = s_387[1:0];
  assign s_461 = {s_462,s_464};
  assign s_462 = s_304 & s_463;
  assign s_463 = ~s_383;
  assign s_464 = s_304?s_465:s_466;
  assign s_465 = s_384[2:0];
  assign s_466 = s_305[2:0];
  assign s_467 = {s_468,s_470};
  assign s_468 = s_119 & s_469;
  assign s_469 = ~s_301;
  assign s_470 = s_119?s_471:s_472;
  assign s_471 = s_302[3:0];
  assign s_472 = s_120[3:0];
  dq #(10, 1) dq_s_473 (clk, s_473, s_474);
  assign s_474 = s_475 - s_478;
  assign s_475 = $signed(s_476);
  assign s_476 = s_108?s_477:s_109;
  assign s_477 = -8'd126;
  assign s_478 = -10'd252;
  assign s_479 = s_480 <= s_481;
  assign s_480 = s_116;
  dq #(10, 1) dq_s_481 (clk, s_481, s_474);
  assign s_482 = 1'd1;
  assign s_483 = s_484[0];
  dq #(10, 1) dq_s_484 (clk, s_484, s_485);
  assign s_485 = s_486 - s_114;
  dq #(10, 2) dq_s_486 (clk, s_486, s_475);
  assign s_487 = 5'd25;
  assign s_488 = 51'd16777216;
  assign s_489 = s_490 <= s_97;
  assign s_490 = s_491 | s_496;
  assign s_491 = s_492 + s_494;
  assign s_492 = s_89?s_493:s_93;
  dq #(52, 3) dq_s_493 (clk, s_493, s_91);
  assign s_494 = s_84 << s_495;
  assign s_495 = 5'd25;
  assign s_496 = 49'd281474976710656;
  assign s_497 = 51'd8388608;
  assign s_498 = s_499 <= s_97;
  assign s_499 = s_500 | s_504;
  assign s_500 = s_501 + s_502;
  assign s_501 = s_489?s_490:s_492;
  assign s_502 = s_82 << s_503;
  assign s_503 = 5'd24;
  assign s_504 = 47'd70368744177664;
  assign s_505 = 51'd4194304;
  assign s_506 = s_507 <= s_97;
  assign s_507 = s_508 | s_512;
  assign s_508 = s_509 + s_510;
  assign s_509 = s_498?s_499:s_501;
  assign s_510 = s_80 << s_511;
  assign s_511 = 5'd23;
  assign s_512 = 45'd17592186044416;
  assign s_513 = 51'd2097152;
  assign s_514 = s_515 <= s_97;
  assign s_515 = s_516 | s_520;
  assign s_516 = s_517 + s_518;
  assign s_517 = s_506?s_507:s_509;
  assign s_518 = s_78 << s_519;
  assign s_519 = 5'd22;
  assign s_520 = 43'd4398046511104;
  assign s_521 = 51'd1048576;
  assign s_522 = s_523 <= s_97;
  assign s_523 = s_524 | s_528;
  assign s_524 = s_525 + s_526;
  assign s_525 = s_514?s_515:s_517;
  assign s_526 = s_76 << s_527;
  assign s_527 = 5'd21;
  assign s_528 = 41'd1099511627776;
  assign s_529 = 51'd524288;
  assign s_530 = s_531 <= s_97;
  assign s_531 = s_532 | s_536;
  assign s_532 = s_533 + s_534;
  assign s_533 = s_522?s_523:s_525;
  assign s_534 = s_74 << s_535;
  assign s_535 = 5'd20;
  assign s_536 = 39'd274877906944;
  assign s_537 = 51'd262144;
  assign s_538 = s_539 <= s_97;
  assign s_539 = s_540 | s_544;
  assign s_540 = s_541 + s_542;
  assign s_541 = s_530?s_531:s_533;
  assign s_542 = s_72 << s_543;
  assign s_543 = 5'd19;
  assign s_544 = 37'd68719476736;
  assign s_545 = 51'd131072;
  assign s_546 = s_547 <= s_97;
  assign s_547 = s_548 | s_552;
  assign s_548 = s_549 + s_550;
  assign s_549 = s_538?s_539:s_541;
  assign s_550 = s_70 << s_551;
  assign s_551 = 5'd18;
  assign s_552 = 35'd17179869184;
  assign s_553 = 51'd65536;
  assign s_554 = s_555 <= s_97;
  assign s_555 = s_556 | s_560;
  assign s_556 = s_557 + s_558;
  assign s_557 = s_546?s_547:s_549;
  assign s_558 = s_68 << s_559;
  assign s_559 = 5'd17;
  assign s_560 = 33'd4294967296;
  assign s_561 = 51'd32768;
  assign s_562 = s_563 <= s_97;
  assign s_563 = s_564 | s_568;
  assign s_564 = s_565 + s_566;
  assign s_565 = s_554?s_555:s_557;
  assign s_566 = s_66 << s_567;
  assign s_567 = 5'd16;
  assign s_568 = 31'd1073741824;
  assign s_569 = 51'd16384;
  assign s_570 = s_571 <= s_97;
  assign s_571 = s_572 | s_576;
  assign s_572 = s_573 + s_574;
  assign s_573 = s_562?s_563:s_565;
  assign s_574 = s_64 << s_575;
  assign s_575 = 4'd15;
  assign s_576 = 29'd268435456;
  assign s_577 = 51'd8192;
  assign s_578 = s_579 <= s_97;
  assign s_579 = s_580 | s_584;
  assign s_580 = s_581 + s_582;
  assign s_581 = s_570?s_571:s_573;
  assign s_582 = s_62 << s_583;
  assign s_583 = 4'd14;
  assign s_584 = 27'd67108864;
  assign s_585 = 51'd4096;
  assign s_586 = s_587 <= s_97;
  assign s_587 = s_588 | s_592;
  assign s_588 = s_589 + s_590;
  assign s_589 = s_578?s_579:s_581;
  assign s_590 = s_60 << s_591;
  assign s_591 = 4'd13;
  assign s_592 = 25'd16777216;
  assign s_593 = 51'd2048;
  assign s_594 = s_595 <= s_97;
  assign s_595 = s_596 | s_600;
  assign s_596 = s_597 + s_598;
  assign s_597 = s_586?s_587:s_589;
  assign s_598 = s_58 << s_599;
  assign s_599 = 4'd12;
  assign s_600 = 23'd4194304;
  assign s_601 = 51'd1024;
  assign s_602 = s_603 <= s_97;
  assign s_603 = s_604 | s_608;
  assign s_604 = s_605 + s_606;
  assign s_605 = s_594?s_595:s_597;
  assign s_606 = s_56 << s_607;
  assign s_607 = 4'd11;
  assign s_608 = 21'd1048576;
  assign s_609 = 51'd512;
  assign s_610 = s_611 <= s_97;
  assign s_611 = s_612 | s_616;
  assign s_612 = s_613 + s_614;
  assign s_613 = s_602?s_603:s_605;
  assign s_614 = s_54 << s_615;
  assign s_615 = 4'd10;
  assign s_616 = 19'd262144;
  assign s_617 = 51'd256;
  assign s_618 = s_619 <= s_97;
  assign s_619 = s_620 | s_624;
  assign s_620 = s_621 + s_622;
  assign s_621 = s_610?s_611:s_613;
  assign s_622 = s_52 << s_623;
  assign s_623 = 4'd9;
  assign s_624 = 17'd65536;
  assign s_625 = 51'd128;
  assign s_626 = s_627 <= s_97;
  assign s_627 = s_628 | s_632;
  assign s_628 = s_629 + s_630;
  assign s_629 = s_618?s_619:s_621;
  assign s_630 = s_50 << s_631;
  assign s_631 = 4'd8;
  assign s_632 = 15'd16384;
  assign s_633 = 51'd64;
  assign s_634 = s_635 <= s_97;
  assign s_635 = s_636 | s_640;
  assign s_636 = s_637 + s_638;
  assign s_637 = s_626?s_627:s_629;
  assign s_638 = s_48 << s_639;
  assign s_639 = 3'd7;
  assign s_640 = 13'd4096;
  assign s_641 = 51'd32;
  assign s_642 = s_643 <= s_97;
  assign s_643 = s_644 | s_648;
  assign s_644 = s_645 + s_646;
  assign s_645 = s_634?s_635:s_637;
  assign s_646 = s_46 << s_647;
  assign s_647 = 3'd6;
  assign s_648 = 11'd1024;
  assign s_649 = 51'd16;
  assign s_650 = s_651 <= s_97;
  assign s_651 = s_652 | s_656;
  assign s_652 = s_653 + s_654;
  assign s_653 = s_642?s_643:s_645;
  assign s_654 = s_44 << s_655;
  assign s_655 = 3'd5;
  assign s_656 = 9'd256;
  assign s_657 = 51'd8;
  assign s_658 = s_659 <= s_97;
  assign s_659 = s_660 | s_664;
  assign s_660 = s_661 + s_662;
  assign s_661 = s_650?s_651:s_653;
  assign s_662 = s_42 << s_663;
  assign s_663 = 3'd4;
  assign s_664 = 7'd64;
  assign s_665 = 51'd4;
  assign s_666 = s_667 <= s_97;
  assign s_667 = s_668 | s_672;
  assign s_668 = s_669 + s_670;
  assign s_669 = s_658?s_659:s_661;
  assign s_670 = s_40 << s_671;
  assign s_671 = 2'd3;
  assign s_672 = 5'd16;
  assign s_673 = 51'd2;
  assign s_674 = s_675 <= s_97;
  assign s_675 = s_676 | s_680;
  assign s_676 = s_677 + s_678;
  assign s_677 = s_666?s_667:s_669;
  assign s_678 = s_38 << s_679;
  assign s_679 = 2'd2;
  assign s_680 = 3'd4;
  assign s_681 = 51'd1;
  assign s_682 = s_683 <= s_97;
  assign s_683 = s_684 | s_688;
  assign s_684 = s_685 + s_686;
  assign s_685 = s_674?s_675:s_677;
  assign s_686 = s_36 << s_687;
  assign s_687 = 1'd1;
  assign s_688 = 1'd1;
  dq #(10, 1) dq_s_689 (clk, s_689, s_690);
  assign s_690 = s_700?s_691:s_692;
  assign s_691 = 1'd0;
  assign s_692 = s_693 - s_694;
  assign s_693 = -10'd126;
  dq #(10, 1) dq_s_694 (clk, s_694, s_695);
  assign s_695 = $signed(s_696) >>> $signed(s_699);
  assign s_696 = s_483?s_697:s_484;
  assign s_697 = s_484 - s_698;
  assign s_698 = 1'd1;
  assign s_699 = 10'd1;
  assign s_700 = s_692[9];
  dq #(10, 1) dq_s_701 (clk, s_701, s_702);
  assign s_702 = s_1064?s_703:s_1058;
  dq #(6, 1) dq_s_703 (clk, s_703, s_704);
  assign s_704 = {s_705,s_1052};
  assign s_705 = s_706 & s_886;
  assign s_706 = s_707[4];
  assign s_707 = {s_708,s_880};
  assign s_708 = s_709 & s_802;
  assign s_709 = s_710[3];
  assign s_710 = {s_711,s_796};
  assign s_711 = s_712 & s_762;
  assign s_712 = s_713[2];
  assign s_713 = {s_714,s_756};
  assign s_714 = s_715 & s_744;
  assign s_715 = s_716[1];
  assign s_716 = {s_717,s_740};
  assign s_717 = s_718 & s_738;
  assign s_718 = ~s_719;
  assign s_719 = s_720[1];
  assign s_720 = s_721[3:2];
  assign s_721 = s_722[7:4];
  assign s_722 = s_723[15:8];
  assign s_723 = s_724[31:16];
  assign s_724 = {s_725,s_737};
  assign s_725 = {s_726,s_736};
  assign s_726 = {s_727,s_735};
  assign s_727 = {s_728,s_734};
  assign s_728 = {s_729,s_733};
  assign s_729 = {s_730,s_732};
  assign s_730 = {s_30,s_731};
  assign s_731 = 1'd1;
  assign s_732 = 1'd1;
  assign s_733 = 1'd1;
  assign s_734 = 1'd1;
  assign s_735 = 1'd1;
  assign s_736 = 1'd1;
  assign s_737 = 1'd1;
  assign s_738 = ~s_739;
  assign s_739 = s_720[0];
  assign s_740 = s_741 & s_743;
  assign s_741 = ~s_742;
  assign s_742 = s_720[1];
  assign s_743 = s_720[0];
  assign s_744 = s_745[1];
  assign s_745 = {s_746,s_752};
  assign s_746 = s_747 & s_750;
  assign s_747 = ~s_748;
  assign s_748 = s_749[1];
  assign s_749 = s_721[1:0];
  assign s_750 = ~s_751;
  assign s_751 = s_749[0];
  assign s_752 = s_753 & s_755;
  assign s_753 = ~s_754;
  assign s_754 = s_749[1];
  assign s_755 = s_749[0];
  assign s_756 = {s_757,s_759};
  assign s_757 = s_715 & s_758;
  assign s_758 = ~s_744;
  assign s_759 = s_715?s_760:s_761;
  assign s_760 = s_745[0:0];
  assign s_761 = s_716[0:0];
  assign s_762 = s_763[2];
  assign s_763 = {s_764,s_790};
  assign s_764 = s_765 & s_778;
  assign s_765 = s_766[1];
  assign s_766 = {s_767,s_774};
  assign s_767 = s_768 & s_772;
  assign s_768 = ~s_769;
  assign s_769 = s_770[1];
  assign s_770 = s_771[3:2];
  assign s_771 = s_722[3:0];
  assign s_772 = ~s_773;
  assign s_773 = s_770[0];
  assign s_774 = s_775 & s_777;
  assign s_775 = ~s_776;
  assign s_776 = s_770[1];
  assign s_777 = s_770[0];
  assign s_778 = s_779[1];
  assign s_779 = {s_780,s_786};
  assign s_780 = s_781 & s_784;
  assign s_781 = ~s_782;
  assign s_782 = s_783[1];
  assign s_783 = s_771[1:0];
  assign s_784 = ~s_785;
  assign s_785 = s_783[0];
  assign s_786 = s_787 & s_789;
  assign s_787 = ~s_788;
  assign s_788 = s_783[1];
  assign s_789 = s_783[0];
  assign s_790 = {s_791,s_793};
  assign s_791 = s_765 & s_792;
  assign s_792 = ~s_778;
  assign s_793 = s_765?s_794:s_795;
  assign s_794 = s_779[0:0];
  assign s_795 = s_766[0:0];
  assign s_796 = {s_797,s_799};
  assign s_797 = s_712 & s_798;
  assign s_798 = ~s_762;
  assign s_799 = s_712?s_800:s_801;
  assign s_800 = s_763[1:0];
  assign s_801 = s_713[1:0];
  assign s_802 = s_803[3];
  assign s_803 = {s_804,s_874};
  assign s_804 = s_805 & s_840;
  assign s_805 = s_806[2];
  assign s_806 = {s_807,s_834};
  assign s_807 = s_808 & s_822;
  assign s_808 = s_809[1];
  assign s_809 = {s_810,s_818};
  assign s_810 = s_811 & s_816;
  assign s_811 = ~s_812;
  assign s_812 = s_813[1];
  assign s_813 = s_814[3:2];
  assign s_814 = s_815[7:4];
  assign s_815 = s_723[7:0];
  assign s_816 = ~s_817;
  assign s_817 = s_813[0];
  assign s_818 = s_819 & s_821;
  assign s_819 = ~s_820;
  assign s_820 = s_813[1];
  assign s_821 = s_813[0];
  assign s_822 = s_823[1];
  assign s_823 = {s_824,s_830};
  assign s_824 = s_825 & s_828;
  assign s_825 = ~s_826;
  assign s_826 = s_827[1];
  assign s_827 = s_814[1:0];
  assign s_828 = ~s_829;
  assign s_829 = s_827[0];
  assign s_830 = s_831 & s_833;
  assign s_831 = ~s_832;
  assign s_832 = s_827[1];
  assign s_833 = s_827[0];
  assign s_834 = {s_835,s_837};
  assign s_835 = s_808 & s_836;
  assign s_836 = ~s_822;
  assign s_837 = s_808?s_838:s_839;
  assign s_838 = s_823[0:0];
  assign s_839 = s_809[0:0];
  assign s_840 = s_841[2];
  assign s_841 = {s_842,s_868};
  assign s_842 = s_843 & s_856;
  assign s_843 = s_844[1];
  assign s_844 = {s_845,s_852};
  assign s_845 = s_846 & s_850;
  assign s_846 = ~s_847;
  assign s_847 = s_848[1];
  assign s_848 = s_849[3:2];
  assign s_849 = s_815[3:0];
  assign s_850 = ~s_851;
  assign s_851 = s_848[0];
  assign s_852 = s_853 & s_855;
  assign s_853 = ~s_854;
  assign s_854 = s_848[1];
  assign s_855 = s_848[0];
  assign s_856 = s_857[1];
  assign s_857 = {s_858,s_864};
  assign s_858 = s_859 & s_862;
  assign s_859 = ~s_860;
  assign s_860 = s_861[1];
  assign s_861 = s_849[1:0];
  assign s_862 = ~s_863;
  assign s_863 = s_861[0];
  assign s_864 = s_865 & s_867;
  assign s_865 = ~s_866;
  assign s_866 = s_861[1];
  assign s_867 = s_861[0];
  assign s_868 = {s_869,s_871};
  assign s_869 = s_843 & s_870;
  assign s_870 = ~s_856;
  assign s_871 = s_843?s_872:s_873;
  assign s_872 = s_857[0:0];
  assign s_873 = s_844[0:0];
  assign s_874 = {s_875,s_877};
  assign s_875 = s_805 & s_876;
  assign s_876 = ~s_840;
  assign s_877 = s_805?s_878:s_879;
  assign s_878 = s_841[1:0];
  assign s_879 = s_806[1:0];
  assign s_880 = {s_881,s_883};
  assign s_881 = s_709 & s_882;
  assign s_882 = ~s_802;
  assign s_883 = s_709?s_884:s_885;
  assign s_884 = s_803[2:0];
  assign s_885 = s_710[2:0];
  assign s_886 = s_887[4];
  assign s_887 = {s_888,s_1046};
  assign s_888 = s_889 & s_968;
  assign s_889 = s_890[3];
  assign s_890 = {s_891,s_962};
  assign s_891 = s_892 & s_928;
  assign s_892 = s_893[2];
  assign s_893 = {s_894,s_922};
  assign s_894 = s_895 & s_910;
  assign s_895 = s_896[1];
  assign s_896 = {s_897,s_906};
  assign s_897 = s_898 & s_904;
  assign s_898 = ~s_899;
  assign s_899 = s_900[1];
  assign s_900 = s_901[3:2];
  assign s_901 = s_902[7:4];
  assign s_902 = s_903[15:8];
  assign s_903 = s_724[15:0];
  assign s_904 = ~s_905;
  assign s_905 = s_900[0];
  assign s_906 = s_907 & s_909;
  assign s_907 = ~s_908;
  assign s_908 = s_900[1];
  assign s_909 = s_900[0];
  assign s_910 = s_911[1];
  assign s_911 = {s_912,s_918};
  assign s_912 = s_913 & s_916;
  assign s_913 = ~s_914;
  assign s_914 = s_915[1];
  assign s_915 = s_901[1:0];
  assign s_916 = ~s_917;
  assign s_917 = s_915[0];
  assign s_918 = s_919 & s_921;
  assign s_919 = ~s_920;
  assign s_920 = s_915[1];
  assign s_921 = s_915[0];
  assign s_922 = {s_923,s_925};
  assign s_923 = s_895 & s_924;
  assign s_924 = ~s_910;
  assign s_925 = s_895?s_926:s_927;
  assign s_926 = s_911[0:0];
  assign s_927 = s_896[0:0];
  assign s_928 = s_929[2];
  assign s_929 = {s_930,s_956};
  assign s_930 = s_931 & s_944;
  assign s_931 = s_932[1];
  assign s_932 = {s_933,s_940};
  assign s_933 = s_934 & s_938;
  assign s_934 = ~s_935;
  assign s_935 = s_936[1];
  assign s_936 = s_937[3:2];
  assign s_937 = s_902[3:0];
  assign s_938 = ~s_939;
  assign s_939 = s_936[0];
  assign s_940 = s_941 & s_943;
  assign s_941 = ~s_942;
  assign s_942 = s_936[1];
  assign s_943 = s_936[0];
  assign s_944 = s_945[1];
  assign s_945 = {s_946,s_952};
  assign s_946 = s_947 & s_950;
  assign s_947 = ~s_948;
  assign s_948 = s_949[1];
  assign s_949 = s_937[1:0];
  assign s_950 = ~s_951;
  assign s_951 = s_949[0];
  assign s_952 = s_953 & s_955;
  assign s_953 = ~s_954;
  assign s_954 = s_949[1];
  assign s_955 = s_949[0];
  assign s_956 = {s_957,s_959};
  assign s_957 = s_931 & s_958;
  assign s_958 = ~s_944;
  assign s_959 = s_931?s_960:s_961;
  assign s_960 = s_945[0:0];
  assign s_961 = s_932[0:0];
  assign s_962 = {s_963,s_965};
  assign s_963 = s_892 & s_964;
  assign s_964 = ~s_928;
  assign s_965 = s_892?s_966:s_967;
  assign s_966 = s_929[1:0];
  assign s_967 = s_893[1:0];
  assign s_968 = s_969[3];
  assign s_969 = {s_970,s_1040};
  assign s_970 = s_971 & s_1006;
  assign s_971 = s_972[2];
  assign s_972 = {s_973,s_1000};
  assign s_973 = s_974 & s_988;
  assign s_974 = s_975[1];
  assign s_975 = {s_976,s_984};
  assign s_976 = s_977 & s_982;
  assign s_977 = ~s_978;
  assign s_978 = s_979[1];
  assign s_979 = s_980[3:2];
  assign s_980 = s_981[7:4];
  assign s_981 = s_903[7:0];
  assign s_982 = ~s_983;
  assign s_983 = s_979[0];
  assign s_984 = s_985 & s_987;
  assign s_985 = ~s_986;
  assign s_986 = s_979[1];
  assign s_987 = s_979[0];
  assign s_988 = s_989[1];
  assign s_989 = {s_990,s_996};
  assign s_990 = s_991 & s_994;
  assign s_991 = ~s_992;
  assign s_992 = s_993[1];
  assign s_993 = s_980[1:0];
  assign s_994 = ~s_995;
  assign s_995 = s_993[0];
  assign s_996 = s_997 & s_999;
  assign s_997 = ~s_998;
  assign s_998 = s_993[1];
  assign s_999 = s_993[0];
  assign s_1000 = {s_1001,s_1003};
  assign s_1001 = s_974 & s_1002;
  assign s_1002 = ~s_988;
  assign s_1003 = s_974?s_1004:s_1005;
  assign s_1004 = s_989[0:0];
  assign s_1005 = s_975[0:0];
  assign s_1006 = s_1007[2];
  assign s_1007 = {s_1008,s_1034};
  assign s_1008 = s_1009 & s_1022;
  assign s_1009 = s_1010[1];
  assign s_1010 = {s_1011,s_1018};
  assign s_1011 = s_1012 & s_1016;
  assign s_1012 = ~s_1013;
  assign s_1013 = s_1014[1];
  assign s_1014 = s_1015[3:2];
  assign s_1015 = s_981[3:0];
  assign s_1016 = ~s_1017;
  assign s_1017 = s_1014[0];
  assign s_1018 = s_1019 & s_1021;
  assign s_1019 = ~s_1020;
  assign s_1020 = s_1014[1];
  assign s_1021 = s_1014[0];
  assign s_1022 = s_1023[1];
  assign s_1023 = {s_1024,s_1030};
  assign s_1024 = s_1025 & s_1028;
  assign s_1025 = ~s_1026;
  assign s_1026 = s_1027[1];
  assign s_1027 = s_1015[1:0];
  assign s_1028 = ~s_1029;
  assign s_1029 = s_1027[0];
  assign s_1030 = s_1031 & s_1033;
  assign s_1031 = ~s_1032;
  assign s_1032 = s_1027[1];
  assign s_1033 = s_1027[0];
  assign s_1034 = {s_1035,s_1037};
  assign s_1035 = s_1009 & s_1036;
  assign s_1036 = ~s_1022;
  assign s_1037 = s_1009?s_1038:s_1039;
  assign s_1038 = s_1023[0:0];
  assign s_1039 = s_1010[0:0];
  assign s_1040 = {s_1041,s_1043};
  assign s_1041 = s_971 & s_1042;
  assign s_1042 = ~s_1006;
  assign s_1043 = s_971?s_1044:s_1045;
  assign s_1044 = s_1007[1:0];
  assign s_1045 = s_972[1:0];
  assign s_1046 = {s_1047,s_1049};
  assign s_1047 = s_889 & s_1048;
  assign s_1048 = ~s_968;
  assign s_1049 = s_889?s_1050:s_1051;
  assign s_1050 = s_969[2:0];
  assign s_1051 = s_890[2:0];
  assign s_1052 = {s_1053,s_1055};
  assign s_1053 = s_706 & s_1054;
  assign s_1054 = ~s_886;
  assign s_1055 = s_706?s_1056:s_1057;
  assign s_1056 = s_887[3:0];
  assign s_1057 = s_707[3:0];
  dq #(10, 1) dq_s_1058 (clk, s_1058, s_1059);
  assign s_1059 = s_1060 - s_1063;
  dq #(10, 1) dq_s_1060 (clk, s_1060, s_1061);
  assign s_1061 = s_1062 + s_689;
  dq #(10, 1) dq_s_1062 (clk, s_1062, s_694);
  assign s_1063 = -10'd126;
  assign s_1064 = s_1065 <= s_1066;
  assign s_1065 = s_703;
  dq #(10, 1) dq_s_1066 (clk, s_1066, s_1059);
  assign s_1067 = 1'd1;
  assign s_1068 = s_1069 & s_1070;
  assign s_1069 = s_27[0];
  assign s_1070 = s_1071 | s_1075;
  dq #(1, 9) dq_s_1071 (clk, s_1071, s_1072);
  assign s_1072 = s_1073 | s_1074;
  assign s_1073 = 1'd1;
  assign s_1074 = 1'd0;
  assign s_1075 = s_26[0];
  assign s_1076 = s_23[23:0];
  assign s_1077 = s_23[24];
  assign s_1078 = {s_1079,s_1089};
  assign s_1079 = {s_1080,s_1081};
  dq #(1, 10) dq_s_1080 (clk, s_1080, s_3);
  assign s_1081 = s_1082 + s_1088;
  assign s_1082 = s_1083[7:0];
  dq #(10, 1) dq_s_1083 (clk, s_1083, s_1084);
  assign s_1084 = s_1085 + s_1077;
  dq #(10, 1) dq_s_1085 (clk, s_1085, s_1086);
  assign s_1086 = s_1087 - s_701;
  dq #(10, 2) dq_s_1087 (clk, s_1087, s_1060);
  assign s_1088 = 7'd127;
  assign s_1089 = s_20[22:0];
  assign s_1090 = s_1091 & s_1093;
  assign s_1091 = s_1082 == s_1092;
  assign s_1092 = -8'd126;
  assign s_1093 = ~s_1094;
  assign s_1094 = s_20[23];
  assign s_1095 = s_20 == s_1096;
  assign s_1096 = 24'd0;
  dq #(1, 10) dq_s_1097 (clk, s_1097, s_1098);
  assign s_1098 = s_1099 & s_1101;
  assign s_1099 = s_109 == s_1100;
  assign s_1100 = 8'd128;
  assign s_1101 = s_113 == s_1102;
  assign s_1102 = 23'd0;
  assign s_1103 = s_1104 | s_1110;
  dq #(1, 10) dq_s_1104 (clk, s_1104, s_1105);
  assign s_1105 = s_1106 & s_1108;
  assign s_1106 = s_109 == s_1107;
  assign s_1107 = 8'd128;
  assign s_1108 = s_113 != s_1109;
  assign s_1109 = 23'd0;
  assign s_1110 = s_1111 & s_1112;
  dq #(1, 10) dq_s_1111 (clk, s_1111, s_3);
  assign s_1112 = s_20 != s_1113;
  assign s_1113 = 1'd0;
  assign sqrt_z = s_0;
endmodule
