module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module lz(clk, a, msb, lsb, msbs_are_zero, lsbs_are_zero, z);
  input clk;
  input [2:0] a;
  output [1:0] msb;
  output [1:0] lsb;
  output [0:0] msbs_are_zero;
  output [0:0] lsbs_are_zero;
  output [2:0] z;
  wire [2:0] s_0;
  wire [0:0] s_1;
  wire [3:0] s_2;
  wire [1:0] s_3;
  wire [1:0] s_4;
  wire [0:0] s_5;
  wire [0:0] s_6;
  wire [0:0] s_7;
  wire [0:0] s_8;
  wire [0:0] s_9;
  wire [0:0] s_10;
  wire [0:0] s_11;
  wire [0:0] s_12;
  wire [0:0] s_13;
  wire [1:0] s_14;
  wire [0:0] s_15;
  wire [0:0] s_16;
  wire [0:0] s_17;
  wire [0:0] s_18;
  wire [0:0] s_19;
  wire [0:0] s_20;
  wire [0:0] s_21;
  wire [0:0] s_22;
  wire [0:0] s_23;
  wire [1:0] s_24;
  wire [0:0] s_25;
  wire [0:0] s_26;
  wire [0:0] s_27;
  wire [0:0] s_28;
  wire [0:0] s_29;
  wire [0:0] s_30;
  wire [0:0] s_31;
  wire [0:0] s_32;
  wire [1:0] s_33;
  wire [2:0] s_34;

  assign s_0 = a;
  assign s_1 = 1'd1;
  assign s_2 = {s_0,s_1};
  assign s_3 = s_2[3:2];
  assign s_4 = s_2[1:0];
  assign s_5 = s_4[1];
  assign s_6 = ~s_5;
  assign s_7 = s_4[0];
  assign s_8 = ~s_7;
  assign s_9 = s_6 & s_8;
  assign s_10 = s_4[1];
  assign s_11 = ~s_10;
  assign s_12 = s_4[0];
  assign s_13 = s_11 & s_12;
  assign s_14 = {s_9,s_13};
  assign s_15 = s_3[1];
  assign s_16 = ~s_15;
  assign s_17 = s_3[0];
  assign s_18 = ~s_17;
  assign s_19 = s_16 & s_18;
  assign s_20 = s_3[1];
  assign s_21 = ~s_20;
  assign s_22 = s_3[0];
  assign s_23 = s_21 & s_22;
  assign s_24 = {s_19,s_23};
  assign s_25 = s_14[1];
  assign s_26 = s_24[1];
  assign s_27 = s_14[0:0];
  assign s_28 = s_24[0:0];
  assign s_29 = s_26 & s_25;
  assign s_30 = ~s_25;
  assign s_31 = s_26 & s_30;
  assign s_32 = s_26?s_27:s_28;
  assign s_33 = {s_31,s_32};
  assign s_34 = {s_29,s_33};
  assign msb = s_3;
  assign lsb = s_4;
  assign msbs_are_zero = s_26;
  assign lsbs_are_zero = s_25;
  assign z = s_34;
endmodule
