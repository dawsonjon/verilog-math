module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module double_div(clk, double_div_a, double_div_b, double_div_z);
  input clk;
  input [63:0] double_div_a;
  input [63:0] double_div_b;
  output [63:0] double_div_z;
  wire [63:0] s_0;
  wire [63:0] s_1;
  wire [63:0] s_2;
  wire [0:0] s_3;
  wire [0:0] s_4;
  wire [63:0] s_5;
  wire [0:0] s_6;
  wire [63:0] s_7;
  wire [62:0] s_8;
  wire [63:0] s_9;
  wire [63:0] s_10;
  wire [63:0] s_11;
  wire [62:0] s_12;
  wire [63:0] s_13;
  wire [63:0] s_14;
  wire [63:0] s_15;
  wire [62:0] s_16;
  wire [63:0] s_17;
  wire [63:0] s_18;
  wire [11:0] s_19;
  wire [11:0] s_20;
  wire [10:0] s_21;
  wire [51:0] s_22;
  wire [52:0] s_23;
  wire [0:0] s_24;
  wire [52:0] s_25;
  wire [52:0] s_26;
  wire [52:0] s_27;
  wire [53:0] s_28;
  wire [53:0] s_29;
  wire [53:0] s_30;
  wire [53:0] s_31;
  wire [52:0] s_32;
  wire [55:0] s_33;
  wire [55:0] s_34;
  wire [55:0] s_35;
  wire [55:0] s_36;
  wire [55:0] s_37;
  wire [55:0] s_38;
  wire [55:0] s_39;
  wire [55:0] s_40;
  wire [55:0] s_41;
  wire [55:0] s_42;
  wire [55:0] s_43;
  wire [55:0] s_44;
  wire [55:0] s_45;
  wire [55:0] s_46;
  wire [55:0] s_47;
  wire [55:0] s_48;
  wire [55:0] s_49;
  wire [55:0] s_50;
  wire [55:0] s_51;
  wire [55:0] s_52;
  wire [55:0] s_53;
  wire [55:0] s_54;
  wire [55:0] s_55;
  wire [55:0] s_56;
  wire [55:0] s_57;
  wire [55:0] s_58;
  wire [55:0] s_59;
  wire [55:0] s_60;
  wire [55:0] s_61;
  wire [55:0] s_62;
  wire [55:0] s_63;
  wire [55:0] s_64;
  wire [55:0] s_65;
  wire [55:0] s_66;
  wire [55:0] s_67;
  wire [55:0] s_68;
  wire [55:0] s_69;
  wire [55:0] s_70;
  wire [55:0] s_71;
  wire [55:0] s_72;
  wire [55:0] s_73;
  wire [55:0] s_74;
  wire [55:0] s_75;
  wire [55:0] s_76;
  wire [55:0] s_77;
  wire [55:0] s_78;
  wire [55:0] s_79;
  wire [55:0] s_80;
  wire [55:0] s_81;
  wire [55:0] s_82;
  wire [55:0] s_83;
  wire [55:0] s_84;
  wire [55:0] s_85;
  wire [55:0] s_86;
  wire [55:0] s_87;
  wire [55:0] s_88;
  wire [55:0] s_89;
  wire [55:0] s_90;
  wire [55:0] s_91;
  wire [55:0] s_92;
  wire [55:0] s_93;
  wire [55:0] s_94;
  wire [55:0] s_95;
  wire [55:0] s_96;
  wire [55:0] s_97;
  wire [55:0] s_98;
  wire [55:0] s_99;
  wire [55:0] s_100;
  wire [55:0] s_101;
  wire [55:0] s_102;
  wire [55:0] s_103;
  wire [55:0] s_104;
  wire [55:0] s_105;
  wire [55:0] s_106;
  wire [55:0] s_107;
  wire [55:0] s_108;
  wire [55:0] s_109;
  wire [55:0] s_110;
  wire [55:0] s_111;
  wire [55:0] s_112;
  wire [55:0] s_113;
  wire [55:0] s_114;
  wire [55:0] s_115;
  wire [55:0] s_116;
  wire [55:0] s_117;
  wire [55:0] s_118;
  wire [55:0] s_119;
  wire [55:0] s_120;
  wire [55:0] s_121;
  wire [55:0] s_122;
  wire [55:0] s_123;
  wire [55:0] s_124;
  wire [55:0] s_125;
  wire [55:0] s_126;
  wire [55:0] s_127;
  wire [55:0] s_128;
  wire [55:0] s_129;
  wire [55:0] s_130;
  wire [55:0] s_131;
  wire [55:0] s_132;
  wire [55:0] s_133;
  wire [55:0] s_134;
  wire [55:0] s_135;
  wire [55:0] s_136;
  wire [55:0] s_137;
  wire [55:0] s_138;
  wire [55:0] s_139;
  wire [55:0] s_140;
  wire [55:0] s_141;
  wire [55:0] s_142;
  wire [55:0] s_143;
  wire [55:0] s_144;
  wire [55:0] s_145;
  wire [55:0] s_146;
  wire [55:0] s_147;
  wire [55:0] s_148;
  wire [55:0] s_149;
  wire [55:0] s_150;
  wire [55:0] s_151;
  wire [55:0] s_152;
  wire [55:0] s_153;
  wire [55:0] s_154;
  wire [55:0] s_155;
  wire [55:0] s_156;
  wire [55:0] s_157;
  wire [55:0] s_158;
  wire [55:0] s_159;
  wire [55:0] s_160;
  wire [55:0] s_161;
  wire [55:0] s_162;
  wire [55:0] s_163;
  wire [55:0] s_164;
  wire [55:0] s_165;
  wire [55:0] s_166;
  wire [55:0] s_167;
  wire [55:0] s_168;
  wire [55:0] s_169;
  wire [55:0] s_170;
  wire [55:0] s_171;
  wire [55:0] s_172;
  wire [55:0] s_173;
  wire [55:0] s_174;
  wire [55:0] s_175;
  wire [55:0] s_176;
  wire [55:0] s_177;
  wire [55:0] s_178;
  wire [55:0] s_179;
  wire [55:0] s_180;
  wire [55:0] s_181;
  wire [55:0] s_182;
  wire [55:0] s_183;
  wire [55:0] s_184;
  wire [55:0] s_185;
  wire [55:0] s_186;
  wire [55:0] s_187;
  wire [55:0] s_188;
  wire [55:0] s_189;
  wire [55:0] s_190;
  wire [55:0] s_191;
  wire [55:0] s_192;
  wire [55:0] s_193;
  wire [55:0] s_194;
  wire [55:0] s_195;
  wire [55:0] s_196;
  wire [55:0] s_197;
  wire [55:0] s_198;
  wire [55:0] s_199;
  wire [55:0] s_200;
  wire [55:0] s_201;
  wire [55:0] s_202;
  wire [55:0] s_203;
  wire [55:0] s_204;
  wire [55:0] s_205;
  wire [55:0] s_206;
  wire [55:0] s_207;
  wire [55:0] s_208;
  wire [0:0] s_209;
  wire [55:0] s_210;
  wire [55:0] s_211;
  wire [0:0] s_212;
  wire [0:0] s_213;
  wire [56:0] s_214;
  wire [56:0] s_215;
  wire [55:0] s_216;
  wire [55:0] s_217;
  wire [52:0] s_218;
  wire [52:0] s_219;
  wire [52:0] s_220;
  wire [52:0] s_221;
  wire [0:0] s_222;
  wire [0:0] s_223;
  wire [0:0] s_224;
  wire [0:0] s_225;
  wire [10:0] s_226;
  wire [10:0] s_227;
  wire [9:0] s_228;
  wire [10:0] s_229;
  wire [51:0] s_230;
  wire [12:0] s_231;
  wire [12:0] s_232;
  wire [6:0] s_233;
  wire [6:0] s_234;
  wire [0:0] s_235;
  wire [0:0] s_236;
  wire [5:0] s_237;
  wire [0:0] s_238;
  wire [0:0] s_239;
  wire [4:0] s_240;
  wire [0:0] s_241;
  wire [0:0] s_242;
  wire [3:0] s_243;
  wire [0:0] s_244;
  wire [0:0] s_245;
  wire [2:0] s_246;
  wire [0:0] s_247;
  wire [0:0] s_248;
  wire [1:0] s_249;
  wire [0:0] s_250;
  wire [0:0] s_251;
  wire [0:0] s_252;
  wire [1:0] s_253;
  wire [3:0] s_254;
  wire [7:0] s_255;
  wire [15:0] s_256;
  wire [31:0] s_257;
  wire [63:0] s_258;
  wire [62:0] s_259;
  wire [61:0] s_260;
  wire [60:0] s_261;
  wire [59:0] s_262;
  wire [58:0] s_263;
  wire [57:0] s_264;
  wire [56:0] s_265;
  wire [55:0] s_266;
  wire [54:0] s_267;
  wire [53:0] s_268;
  wire [0:0] s_269;
  wire [0:0] s_270;
  wire [0:0] s_271;
  wire [0:0] s_272;
  wire [0:0] s_273;
  wire [0:0] s_274;
  wire [0:0] s_275;
  wire [0:0] s_276;
  wire [0:0] s_277;
  wire [0:0] s_278;
  wire [0:0] s_279;
  wire [0:0] s_280;
  wire [0:0] s_281;
  wire [0:0] s_282;
  wire [0:0] s_283;
  wire [0:0] s_284;
  wire [0:0] s_285;
  wire [0:0] s_286;
  wire [1:0] s_287;
  wire [0:0] s_288;
  wire [0:0] s_289;
  wire [0:0] s_290;
  wire [1:0] s_291;
  wire [0:0] s_292;
  wire [0:0] s_293;
  wire [0:0] s_294;
  wire [0:0] s_295;
  wire [0:0] s_296;
  wire [0:0] s_297;
  wire [1:0] s_298;
  wire [0:0] s_299;
  wire [0:0] s_300;
  wire [0:0] s_301;
  wire [0:0] s_302;
  wire [0:0] s_303;
  wire [0:0] s_304;
  wire [2:0] s_305;
  wire [0:0] s_306;
  wire [0:0] s_307;
  wire [1:0] s_308;
  wire [0:0] s_309;
  wire [0:0] s_310;
  wire [0:0] s_311;
  wire [1:0] s_312;
  wire [3:0] s_313;
  wire [0:0] s_314;
  wire [0:0] s_315;
  wire [0:0] s_316;
  wire [0:0] s_317;
  wire [0:0] s_318;
  wire [0:0] s_319;
  wire [0:0] s_320;
  wire [1:0] s_321;
  wire [0:0] s_322;
  wire [0:0] s_323;
  wire [0:0] s_324;
  wire [1:0] s_325;
  wire [0:0] s_326;
  wire [0:0] s_327;
  wire [0:0] s_328;
  wire [0:0] s_329;
  wire [0:0] s_330;
  wire [0:0] s_331;
  wire [1:0] s_332;
  wire [0:0] s_333;
  wire [0:0] s_334;
  wire [0:0] s_335;
  wire [0:0] s_336;
  wire [0:0] s_337;
  wire [2:0] s_338;
  wire [0:0] s_339;
  wire [0:0] s_340;
  wire [1:0] s_341;
  wire [1:0] s_342;
  wire [1:0] s_343;
  wire [0:0] s_344;
  wire [3:0] s_345;
  wire [0:0] s_346;
  wire [0:0] s_347;
  wire [2:0] s_348;
  wire [0:0] s_349;
  wire [0:0] s_350;
  wire [1:0] s_351;
  wire [0:0] s_352;
  wire [0:0] s_353;
  wire [0:0] s_354;
  wire [1:0] s_355;
  wire [3:0] s_356;
  wire [7:0] s_357;
  wire [0:0] s_358;
  wire [0:0] s_359;
  wire [0:0] s_360;
  wire [0:0] s_361;
  wire [0:0] s_362;
  wire [0:0] s_363;
  wire [0:0] s_364;
  wire [1:0] s_365;
  wire [0:0] s_366;
  wire [0:0] s_367;
  wire [0:0] s_368;
  wire [1:0] s_369;
  wire [0:0] s_370;
  wire [0:0] s_371;
  wire [0:0] s_372;
  wire [0:0] s_373;
  wire [0:0] s_374;
  wire [0:0] s_375;
  wire [1:0] s_376;
  wire [0:0] s_377;
  wire [0:0] s_378;
  wire [0:0] s_379;
  wire [0:0] s_380;
  wire [0:0] s_381;
  wire [0:0] s_382;
  wire [2:0] s_383;
  wire [0:0] s_384;
  wire [0:0] s_385;
  wire [1:0] s_386;
  wire [0:0] s_387;
  wire [0:0] s_388;
  wire [0:0] s_389;
  wire [1:0] s_390;
  wire [3:0] s_391;
  wire [0:0] s_392;
  wire [0:0] s_393;
  wire [0:0] s_394;
  wire [0:0] s_395;
  wire [0:0] s_396;
  wire [0:0] s_397;
  wire [0:0] s_398;
  wire [1:0] s_399;
  wire [0:0] s_400;
  wire [0:0] s_401;
  wire [0:0] s_402;
  wire [1:0] s_403;
  wire [0:0] s_404;
  wire [0:0] s_405;
  wire [0:0] s_406;
  wire [0:0] s_407;
  wire [0:0] s_408;
  wire [0:0] s_409;
  wire [1:0] s_410;
  wire [0:0] s_411;
  wire [0:0] s_412;
  wire [0:0] s_413;
  wire [0:0] s_414;
  wire [0:0] s_415;
  wire [2:0] s_416;
  wire [0:0] s_417;
  wire [0:0] s_418;
  wire [1:0] s_419;
  wire [1:0] s_420;
  wire [1:0] s_421;
  wire [3:0] s_422;
  wire [0:0] s_423;
  wire [0:0] s_424;
  wire [2:0] s_425;
  wire [2:0] s_426;
  wire [2:0] s_427;
  wire [0:0] s_428;
  wire [4:0] s_429;
  wire [0:0] s_430;
  wire [0:0] s_431;
  wire [3:0] s_432;
  wire [0:0] s_433;
  wire [0:0] s_434;
  wire [2:0] s_435;
  wire [0:0] s_436;
  wire [0:0] s_437;
  wire [1:0] s_438;
  wire [0:0] s_439;
  wire [0:0] s_440;
  wire [0:0] s_441;
  wire [1:0] s_442;
  wire [3:0] s_443;
  wire [7:0] s_444;
  wire [15:0] s_445;
  wire [0:0] s_446;
  wire [0:0] s_447;
  wire [0:0] s_448;
  wire [0:0] s_449;
  wire [0:0] s_450;
  wire [0:0] s_451;
  wire [0:0] s_452;
  wire [1:0] s_453;
  wire [0:0] s_454;
  wire [0:0] s_455;
  wire [0:0] s_456;
  wire [1:0] s_457;
  wire [0:0] s_458;
  wire [0:0] s_459;
  wire [0:0] s_460;
  wire [0:0] s_461;
  wire [0:0] s_462;
  wire [0:0] s_463;
  wire [1:0] s_464;
  wire [0:0] s_465;
  wire [0:0] s_466;
  wire [0:0] s_467;
  wire [0:0] s_468;
  wire [0:0] s_469;
  wire [0:0] s_470;
  wire [2:0] s_471;
  wire [0:0] s_472;
  wire [0:0] s_473;
  wire [1:0] s_474;
  wire [0:0] s_475;
  wire [0:0] s_476;
  wire [0:0] s_477;
  wire [1:0] s_478;
  wire [3:0] s_479;
  wire [0:0] s_480;
  wire [0:0] s_481;
  wire [0:0] s_482;
  wire [0:0] s_483;
  wire [0:0] s_484;
  wire [0:0] s_485;
  wire [0:0] s_486;
  wire [1:0] s_487;
  wire [0:0] s_488;
  wire [0:0] s_489;
  wire [0:0] s_490;
  wire [1:0] s_491;
  wire [0:0] s_492;
  wire [0:0] s_493;
  wire [0:0] s_494;
  wire [0:0] s_495;
  wire [0:0] s_496;
  wire [0:0] s_497;
  wire [1:0] s_498;
  wire [0:0] s_499;
  wire [0:0] s_500;
  wire [0:0] s_501;
  wire [0:0] s_502;
  wire [0:0] s_503;
  wire [2:0] s_504;
  wire [0:0] s_505;
  wire [0:0] s_506;
  wire [1:0] s_507;
  wire [1:0] s_508;
  wire [1:0] s_509;
  wire [0:0] s_510;
  wire [3:0] s_511;
  wire [0:0] s_512;
  wire [0:0] s_513;
  wire [2:0] s_514;
  wire [0:0] s_515;
  wire [0:0] s_516;
  wire [1:0] s_517;
  wire [0:0] s_518;
  wire [0:0] s_519;
  wire [0:0] s_520;
  wire [1:0] s_521;
  wire [3:0] s_522;
  wire [7:0] s_523;
  wire [0:0] s_524;
  wire [0:0] s_525;
  wire [0:0] s_526;
  wire [0:0] s_527;
  wire [0:0] s_528;
  wire [0:0] s_529;
  wire [0:0] s_530;
  wire [1:0] s_531;
  wire [0:0] s_532;
  wire [0:0] s_533;
  wire [0:0] s_534;
  wire [1:0] s_535;
  wire [0:0] s_536;
  wire [0:0] s_537;
  wire [0:0] s_538;
  wire [0:0] s_539;
  wire [0:0] s_540;
  wire [0:0] s_541;
  wire [1:0] s_542;
  wire [0:0] s_543;
  wire [0:0] s_544;
  wire [0:0] s_545;
  wire [0:0] s_546;
  wire [0:0] s_547;
  wire [0:0] s_548;
  wire [2:0] s_549;
  wire [0:0] s_550;
  wire [0:0] s_551;
  wire [1:0] s_552;
  wire [0:0] s_553;
  wire [0:0] s_554;
  wire [0:0] s_555;
  wire [1:0] s_556;
  wire [3:0] s_557;
  wire [0:0] s_558;
  wire [0:0] s_559;
  wire [0:0] s_560;
  wire [0:0] s_561;
  wire [0:0] s_562;
  wire [0:0] s_563;
  wire [0:0] s_564;
  wire [1:0] s_565;
  wire [0:0] s_566;
  wire [0:0] s_567;
  wire [0:0] s_568;
  wire [1:0] s_569;
  wire [0:0] s_570;
  wire [0:0] s_571;
  wire [0:0] s_572;
  wire [0:0] s_573;
  wire [0:0] s_574;
  wire [0:0] s_575;
  wire [1:0] s_576;
  wire [0:0] s_577;
  wire [0:0] s_578;
  wire [0:0] s_579;
  wire [0:0] s_580;
  wire [0:0] s_581;
  wire [2:0] s_582;
  wire [0:0] s_583;
  wire [0:0] s_584;
  wire [1:0] s_585;
  wire [1:0] s_586;
  wire [1:0] s_587;
  wire [3:0] s_588;
  wire [0:0] s_589;
  wire [0:0] s_590;
  wire [2:0] s_591;
  wire [2:0] s_592;
  wire [2:0] s_593;
  wire [4:0] s_594;
  wire [0:0] s_595;
  wire [0:0] s_596;
  wire [3:0] s_597;
  wire [3:0] s_598;
  wire [3:0] s_599;
  wire [0:0] s_600;
  wire [5:0] s_601;
  wire [0:0] s_602;
  wire [0:0] s_603;
  wire [4:0] s_604;
  wire [0:0] s_605;
  wire [0:0] s_606;
  wire [3:0] s_607;
  wire [0:0] s_608;
  wire [0:0] s_609;
  wire [2:0] s_610;
  wire [0:0] s_611;
  wire [0:0] s_612;
  wire [1:0] s_613;
  wire [0:0] s_614;
  wire [0:0] s_615;
  wire [0:0] s_616;
  wire [1:0] s_617;
  wire [3:0] s_618;
  wire [7:0] s_619;
  wire [15:0] s_620;
  wire [31:0] s_621;
  wire [0:0] s_622;
  wire [0:0] s_623;
  wire [0:0] s_624;
  wire [0:0] s_625;
  wire [0:0] s_626;
  wire [0:0] s_627;
  wire [0:0] s_628;
  wire [1:0] s_629;
  wire [0:0] s_630;
  wire [0:0] s_631;
  wire [0:0] s_632;
  wire [1:0] s_633;
  wire [0:0] s_634;
  wire [0:0] s_635;
  wire [0:0] s_636;
  wire [0:0] s_637;
  wire [0:0] s_638;
  wire [0:0] s_639;
  wire [1:0] s_640;
  wire [0:0] s_641;
  wire [0:0] s_642;
  wire [0:0] s_643;
  wire [0:0] s_644;
  wire [0:0] s_645;
  wire [0:0] s_646;
  wire [2:0] s_647;
  wire [0:0] s_648;
  wire [0:0] s_649;
  wire [1:0] s_650;
  wire [0:0] s_651;
  wire [0:0] s_652;
  wire [0:0] s_653;
  wire [1:0] s_654;
  wire [3:0] s_655;
  wire [0:0] s_656;
  wire [0:0] s_657;
  wire [0:0] s_658;
  wire [0:0] s_659;
  wire [0:0] s_660;
  wire [0:0] s_661;
  wire [0:0] s_662;
  wire [1:0] s_663;
  wire [0:0] s_664;
  wire [0:0] s_665;
  wire [0:0] s_666;
  wire [1:0] s_667;
  wire [0:0] s_668;
  wire [0:0] s_669;
  wire [0:0] s_670;
  wire [0:0] s_671;
  wire [0:0] s_672;
  wire [0:0] s_673;
  wire [1:0] s_674;
  wire [0:0] s_675;
  wire [0:0] s_676;
  wire [0:0] s_677;
  wire [0:0] s_678;
  wire [0:0] s_679;
  wire [2:0] s_680;
  wire [0:0] s_681;
  wire [0:0] s_682;
  wire [1:0] s_683;
  wire [1:0] s_684;
  wire [1:0] s_685;
  wire [0:0] s_686;
  wire [3:0] s_687;
  wire [0:0] s_688;
  wire [0:0] s_689;
  wire [2:0] s_690;
  wire [0:0] s_691;
  wire [0:0] s_692;
  wire [1:0] s_693;
  wire [0:0] s_694;
  wire [0:0] s_695;
  wire [0:0] s_696;
  wire [1:0] s_697;
  wire [3:0] s_698;
  wire [7:0] s_699;
  wire [0:0] s_700;
  wire [0:0] s_701;
  wire [0:0] s_702;
  wire [0:0] s_703;
  wire [0:0] s_704;
  wire [0:0] s_705;
  wire [0:0] s_706;
  wire [1:0] s_707;
  wire [0:0] s_708;
  wire [0:0] s_709;
  wire [0:0] s_710;
  wire [1:0] s_711;
  wire [0:0] s_712;
  wire [0:0] s_713;
  wire [0:0] s_714;
  wire [0:0] s_715;
  wire [0:0] s_716;
  wire [0:0] s_717;
  wire [1:0] s_718;
  wire [0:0] s_719;
  wire [0:0] s_720;
  wire [0:0] s_721;
  wire [0:0] s_722;
  wire [0:0] s_723;
  wire [0:0] s_724;
  wire [2:0] s_725;
  wire [0:0] s_726;
  wire [0:0] s_727;
  wire [1:0] s_728;
  wire [0:0] s_729;
  wire [0:0] s_730;
  wire [0:0] s_731;
  wire [1:0] s_732;
  wire [3:0] s_733;
  wire [0:0] s_734;
  wire [0:0] s_735;
  wire [0:0] s_736;
  wire [0:0] s_737;
  wire [0:0] s_738;
  wire [0:0] s_739;
  wire [0:0] s_740;
  wire [1:0] s_741;
  wire [0:0] s_742;
  wire [0:0] s_743;
  wire [0:0] s_744;
  wire [1:0] s_745;
  wire [0:0] s_746;
  wire [0:0] s_747;
  wire [0:0] s_748;
  wire [0:0] s_749;
  wire [0:0] s_750;
  wire [0:0] s_751;
  wire [1:0] s_752;
  wire [0:0] s_753;
  wire [0:0] s_754;
  wire [0:0] s_755;
  wire [0:0] s_756;
  wire [0:0] s_757;
  wire [2:0] s_758;
  wire [0:0] s_759;
  wire [0:0] s_760;
  wire [1:0] s_761;
  wire [1:0] s_762;
  wire [1:0] s_763;
  wire [3:0] s_764;
  wire [0:0] s_765;
  wire [0:0] s_766;
  wire [2:0] s_767;
  wire [2:0] s_768;
  wire [2:0] s_769;
  wire [0:0] s_770;
  wire [4:0] s_771;
  wire [0:0] s_772;
  wire [0:0] s_773;
  wire [3:0] s_774;
  wire [0:0] s_775;
  wire [0:0] s_776;
  wire [2:0] s_777;
  wire [0:0] s_778;
  wire [0:0] s_779;
  wire [1:0] s_780;
  wire [0:0] s_781;
  wire [0:0] s_782;
  wire [0:0] s_783;
  wire [1:0] s_784;
  wire [3:0] s_785;
  wire [7:0] s_786;
  wire [15:0] s_787;
  wire [0:0] s_788;
  wire [0:0] s_789;
  wire [0:0] s_790;
  wire [0:0] s_791;
  wire [0:0] s_792;
  wire [0:0] s_793;
  wire [0:0] s_794;
  wire [1:0] s_795;
  wire [0:0] s_796;
  wire [0:0] s_797;
  wire [0:0] s_798;
  wire [1:0] s_799;
  wire [0:0] s_800;
  wire [0:0] s_801;
  wire [0:0] s_802;
  wire [0:0] s_803;
  wire [0:0] s_804;
  wire [0:0] s_805;
  wire [1:0] s_806;
  wire [0:0] s_807;
  wire [0:0] s_808;
  wire [0:0] s_809;
  wire [0:0] s_810;
  wire [0:0] s_811;
  wire [0:0] s_812;
  wire [2:0] s_813;
  wire [0:0] s_814;
  wire [0:0] s_815;
  wire [1:0] s_816;
  wire [0:0] s_817;
  wire [0:0] s_818;
  wire [0:0] s_819;
  wire [1:0] s_820;
  wire [3:0] s_821;
  wire [0:0] s_822;
  wire [0:0] s_823;
  wire [0:0] s_824;
  wire [0:0] s_825;
  wire [0:0] s_826;
  wire [0:0] s_827;
  wire [0:0] s_828;
  wire [1:0] s_829;
  wire [0:0] s_830;
  wire [0:0] s_831;
  wire [0:0] s_832;
  wire [1:0] s_833;
  wire [0:0] s_834;
  wire [0:0] s_835;
  wire [0:0] s_836;
  wire [0:0] s_837;
  wire [0:0] s_838;
  wire [0:0] s_839;
  wire [1:0] s_840;
  wire [0:0] s_841;
  wire [0:0] s_842;
  wire [0:0] s_843;
  wire [0:0] s_844;
  wire [0:0] s_845;
  wire [2:0] s_846;
  wire [0:0] s_847;
  wire [0:0] s_848;
  wire [1:0] s_849;
  wire [1:0] s_850;
  wire [1:0] s_851;
  wire [0:0] s_852;
  wire [3:0] s_853;
  wire [0:0] s_854;
  wire [0:0] s_855;
  wire [2:0] s_856;
  wire [0:0] s_857;
  wire [0:0] s_858;
  wire [1:0] s_859;
  wire [0:0] s_860;
  wire [0:0] s_861;
  wire [0:0] s_862;
  wire [1:0] s_863;
  wire [3:0] s_864;
  wire [7:0] s_865;
  wire [0:0] s_866;
  wire [0:0] s_867;
  wire [0:0] s_868;
  wire [0:0] s_869;
  wire [0:0] s_870;
  wire [0:0] s_871;
  wire [0:0] s_872;
  wire [1:0] s_873;
  wire [0:0] s_874;
  wire [0:0] s_875;
  wire [0:0] s_876;
  wire [1:0] s_877;
  wire [0:0] s_878;
  wire [0:0] s_879;
  wire [0:0] s_880;
  wire [0:0] s_881;
  wire [0:0] s_882;
  wire [0:0] s_883;
  wire [1:0] s_884;
  wire [0:0] s_885;
  wire [0:0] s_886;
  wire [0:0] s_887;
  wire [0:0] s_888;
  wire [0:0] s_889;
  wire [0:0] s_890;
  wire [2:0] s_891;
  wire [0:0] s_892;
  wire [0:0] s_893;
  wire [1:0] s_894;
  wire [0:0] s_895;
  wire [0:0] s_896;
  wire [0:0] s_897;
  wire [1:0] s_898;
  wire [3:0] s_899;
  wire [0:0] s_900;
  wire [0:0] s_901;
  wire [0:0] s_902;
  wire [0:0] s_903;
  wire [0:0] s_904;
  wire [0:0] s_905;
  wire [0:0] s_906;
  wire [1:0] s_907;
  wire [0:0] s_908;
  wire [0:0] s_909;
  wire [0:0] s_910;
  wire [1:0] s_911;
  wire [0:0] s_912;
  wire [0:0] s_913;
  wire [0:0] s_914;
  wire [0:0] s_915;
  wire [0:0] s_916;
  wire [0:0] s_917;
  wire [1:0] s_918;
  wire [0:0] s_919;
  wire [0:0] s_920;
  wire [0:0] s_921;
  wire [0:0] s_922;
  wire [0:0] s_923;
  wire [2:0] s_924;
  wire [0:0] s_925;
  wire [0:0] s_926;
  wire [1:0] s_927;
  wire [1:0] s_928;
  wire [1:0] s_929;
  wire [3:0] s_930;
  wire [0:0] s_931;
  wire [0:0] s_932;
  wire [2:0] s_933;
  wire [2:0] s_934;
  wire [2:0] s_935;
  wire [4:0] s_936;
  wire [0:0] s_937;
  wire [0:0] s_938;
  wire [3:0] s_939;
  wire [3:0] s_940;
  wire [3:0] s_941;
  wire [5:0] s_942;
  wire [0:0] s_943;
  wire [0:0] s_944;
  wire [4:0] s_945;
  wire [4:0] s_946;
  wire [4:0] s_947;
  wire [12:0] s_948;
  wire [12:0] s_949;
  wire [12:0] s_950;
  wire [10:0] s_951;
  wire [10:0] s_952;
  wire [12:0] s_953;
  wire [0:0] s_954;
  wire [12:0] s_955;
  wire [12:0] s_956;
  wire [1:0] s_957;
  wire [55:0] s_958;
  wire [55:0] s_959;
  wire [52:0] s_960;
  wire [52:0] s_961;
  wire [52:0] s_962;
  wire [52:0] s_963;
  wire [0:0] s_964;
  wire [0:0] s_965;
  wire [0:0] s_966;
  wire [0:0] s_967;
  wire [10:0] s_968;
  wire [10:0] s_969;
  wire [9:0] s_970;
  wire [10:0] s_971;
  wire [51:0] s_972;
  wire [12:0] s_973;
  wire [12:0] s_974;
  wire [6:0] s_975;
  wire [6:0] s_976;
  wire [0:0] s_977;
  wire [0:0] s_978;
  wire [5:0] s_979;
  wire [0:0] s_980;
  wire [0:0] s_981;
  wire [4:0] s_982;
  wire [0:0] s_983;
  wire [0:0] s_984;
  wire [3:0] s_985;
  wire [0:0] s_986;
  wire [0:0] s_987;
  wire [2:0] s_988;
  wire [0:0] s_989;
  wire [0:0] s_990;
  wire [1:0] s_991;
  wire [0:0] s_992;
  wire [0:0] s_993;
  wire [0:0] s_994;
  wire [1:0] s_995;
  wire [3:0] s_996;
  wire [7:0] s_997;
  wire [15:0] s_998;
  wire [31:0] s_999;
  wire [63:0] s_1000;
  wire [62:0] s_1001;
  wire [61:0] s_1002;
  wire [60:0] s_1003;
  wire [59:0] s_1004;
  wire [58:0] s_1005;
  wire [57:0] s_1006;
  wire [56:0] s_1007;
  wire [55:0] s_1008;
  wire [54:0] s_1009;
  wire [53:0] s_1010;
  wire [0:0] s_1011;
  wire [0:0] s_1012;
  wire [0:0] s_1013;
  wire [0:0] s_1014;
  wire [0:0] s_1015;
  wire [0:0] s_1016;
  wire [0:0] s_1017;
  wire [0:0] s_1018;
  wire [0:0] s_1019;
  wire [0:0] s_1020;
  wire [0:0] s_1021;
  wire [0:0] s_1022;
  wire [0:0] s_1023;
  wire [0:0] s_1024;
  wire [0:0] s_1025;
  wire [0:0] s_1026;
  wire [0:0] s_1027;
  wire [0:0] s_1028;
  wire [1:0] s_1029;
  wire [0:0] s_1030;
  wire [0:0] s_1031;
  wire [0:0] s_1032;
  wire [1:0] s_1033;
  wire [0:0] s_1034;
  wire [0:0] s_1035;
  wire [0:0] s_1036;
  wire [0:0] s_1037;
  wire [0:0] s_1038;
  wire [0:0] s_1039;
  wire [1:0] s_1040;
  wire [0:0] s_1041;
  wire [0:0] s_1042;
  wire [0:0] s_1043;
  wire [0:0] s_1044;
  wire [0:0] s_1045;
  wire [0:0] s_1046;
  wire [2:0] s_1047;
  wire [0:0] s_1048;
  wire [0:0] s_1049;
  wire [1:0] s_1050;
  wire [0:0] s_1051;
  wire [0:0] s_1052;
  wire [0:0] s_1053;
  wire [1:0] s_1054;
  wire [3:0] s_1055;
  wire [0:0] s_1056;
  wire [0:0] s_1057;
  wire [0:0] s_1058;
  wire [0:0] s_1059;
  wire [0:0] s_1060;
  wire [0:0] s_1061;
  wire [0:0] s_1062;
  wire [1:0] s_1063;
  wire [0:0] s_1064;
  wire [0:0] s_1065;
  wire [0:0] s_1066;
  wire [1:0] s_1067;
  wire [0:0] s_1068;
  wire [0:0] s_1069;
  wire [0:0] s_1070;
  wire [0:0] s_1071;
  wire [0:0] s_1072;
  wire [0:0] s_1073;
  wire [1:0] s_1074;
  wire [0:0] s_1075;
  wire [0:0] s_1076;
  wire [0:0] s_1077;
  wire [0:0] s_1078;
  wire [0:0] s_1079;
  wire [2:0] s_1080;
  wire [0:0] s_1081;
  wire [0:0] s_1082;
  wire [1:0] s_1083;
  wire [1:0] s_1084;
  wire [1:0] s_1085;
  wire [0:0] s_1086;
  wire [3:0] s_1087;
  wire [0:0] s_1088;
  wire [0:0] s_1089;
  wire [2:0] s_1090;
  wire [0:0] s_1091;
  wire [0:0] s_1092;
  wire [1:0] s_1093;
  wire [0:0] s_1094;
  wire [0:0] s_1095;
  wire [0:0] s_1096;
  wire [1:0] s_1097;
  wire [3:0] s_1098;
  wire [7:0] s_1099;
  wire [0:0] s_1100;
  wire [0:0] s_1101;
  wire [0:0] s_1102;
  wire [0:0] s_1103;
  wire [0:0] s_1104;
  wire [0:0] s_1105;
  wire [0:0] s_1106;
  wire [1:0] s_1107;
  wire [0:0] s_1108;
  wire [0:0] s_1109;
  wire [0:0] s_1110;
  wire [1:0] s_1111;
  wire [0:0] s_1112;
  wire [0:0] s_1113;
  wire [0:0] s_1114;
  wire [0:0] s_1115;
  wire [0:0] s_1116;
  wire [0:0] s_1117;
  wire [1:0] s_1118;
  wire [0:0] s_1119;
  wire [0:0] s_1120;
  wire [0:0] s_1121;
  wire [0:0] s_1122;
  wire [0:0] s_1123;
  wire [0:0] s_1124;
  wire [2:0] s_1125;
  wire [0:0] s_1126;
  wire [0:0] s_1127;
  wire [1:0] s_1128;
  wire [0:0] s_1129;
  wire [0:0] s_1130;
  wire [0:0] s_1131;
  wire [1:0] s_1132;
  wire [3:0] s_1133;
  wire [0:0] s_1134;
  wire [0:0] s_1135;
  wire [0:0] s_1136;
  wire [0:0] s_1137;
  wire [0:0] s_1138;
  wire [0:0] s_1139;
  wire [0:0] s_1140;
  wire [1:0] s_1141;
  wire [0:0] s_1142;
  wire [0:0] s_1143;
  wire [0:0] s_1144;
  wire [1:0] s_1145;
  wire [0:0] s_1146;
  wire [0:0] s_1147;
  wire [0:0] s_1148;
  wire [0:0] s_1149;
  wire [0:0] s_1150;
  wire [0:0] s_1151;
  wire [1:0] s_1152;
  wire [0:0] s_1153;
  wire [0:0] s_1154;
  wire [0:0] s_1155;
  wire [0:0] s_1156;
  wire [0:0] s_1157;
  wire [2:0] s_1158;
  wire [0:0] s_1159;
  wire [0:0] s_1160;
  wire [1:0] s_1161;
  wire [1:0] s_1162;
  wire [1:0] s_1163;
  wire [3:0] s_1164;
  wire [0:0] s_1165;
  wire [0:0] s_1166;
  wire [2:0] s_1167;
  wire [2:0] s_1168;
  wire [2:0] s_1169;
  wire [0:0] s_1170;
  wire [4:0] s_1171;
  wire [0:0] s_1172;
  wire [0:0] s_1173;
  wire [3:0] s_1174;
  wire [0:0] s_1175;
  wire [0:0] s_1176;
  wire [2:0] s_1177;
  wire [0:0] s_1178;
  wire [0:0] s_1179;
  wire [1:0] s_1180;
  wire [0:0] s_1181;
  wire [0:0] s_1182;
  wire [0:0] s_1183;
  wire [1:0] s_1184;
  wire [3:0] s_1185;
  wire [7:0] s_1186;
  wire [15:0] s_1187;
  wire [0:0] s_1188;
  wire [0:0] s_1189;
  wire [0:0] s_1190;
  wire [0:0] s_1191;
  wire [0:0] s_1192;
  wire [0:0] s_1193;
  wire [0:0] s_1194;
  wire [1:0] s_1195;
  wire [0:0] s_1196;
  wire [0:0] s_1197;
  wire [0:0] s_1198;
  wire [1:0] s_1199;
  wire [0:0] s_1200;
  wire [0:0] s_1201;
  wire [0:0] s_1202;
  wire [0:0] s_1203;
  wire [0:0] s_1204;
  wire [0:0] s_1205;
  wire [1:0] s_1206;
  wire [0:0] s_1207;
  wire [0:0] s_1208;
  wire [0:0] s_1209;
  wire [0:0] s_1210;
  wire [0:0] s_1211;
  wire [0:0] s_1212;
  wire [2:0] s_1213;
  wire [0:0] s_1214;
  wire [0:0] s_1215;
  wire [1:0] s_1216;
  wire [0:0] s_1217;
  wire [0:0] s_1218;
  wire [0:0] s_1219;
  wire [1:0] s_1220;
  wire [3:0] s_1221;
  wire [0:0] s_1222;
  wire [0:0] s_1223;
  wire [0:0] s_1224;
  wire [0:0] s_1225;
  wire [0:0] s_1226;
  wire [0:0] s_1227;
  wire [0:0] s_1228;
  wire [1:0] s_1229;
  wire [0:0] s_1230;
  wire [0:0] s_1231;
  wire [0:0] s_1232;
  wire [1:0] s_1233;
  wire [0:0] s_1234;
  wire [0:0] s_1235;
  wire [0:0] s_1236;
  wire [0:0] s_1237;
  wire [0:0] s_1238;
  wire [0:0] s_1239;
  wire [1:0] s_1240;
  wire [0:0] s_1241;
  wire [0:0] s_1242;
  wire [0:0] s_1243;
  wire [0:0] s_1244;
  wire [0:0] s_1245;
  wire [2:0] s_1246;
  wire [0:0] s_1247;
  wire [0:0] s_1248;
  wire [1:0] s_1249;
  wire [1:0] s_1250;
  wire [1:0] s_1251;
  wire [0:0] s_1252;
  wire [3:0] s_1253;
  wire [0:0] s_1254;
  wire [0:0] s_1255;
  wire [2:0] s_1256;
  wire [0:0] s_1257;
  wire [0:0] s_1258;
  wire [1:0] s_1259;
  wire [0:0] s_1260;
  wire [0:0] s_1261;
  wire [0:0] s_1262;
  wire [1:0] s_1263;
  wire [3:0] s_1264;
  wire [7:0] s_1265;
  wire [0:0] s_1266;
  wire [0:0] s_1267;
  wire [0:0] s_1268;
  wire [0:0] s_1269;
  wire [0:0] s_1270;
  wire [0:0] s_1271;
  wire [0:0] s_1272;
  wire [1:0] s_1273;
  wire [0:0] s_1274;
  wire [0:0] s_1275;
  wire [0:0] s_1276;
  wire [1:0] s_1277;
  wire [0:0] s_1278;
  wire [0:0] s_1279;
  wire [0:0] s_1280;
  wire [0:0] s_1281;
  wire [0:0] s_1282;
  wire [0:0] s_1283;
  wire [1:0] s_1284;
  wire [0:0] s_1285;
  wire [0:0] s_1286;
  wire [0:0] s_1287;
  wire [0:0] s_1288;
  wire [0:0] s_1289;
  wire [0:0] s_1290;
  wire [2:0] s_1291;
  wire [0:0] s_1292;
  wire [0:0] s_1293;
  wire [1:0] s_1294;
  wire [0:0] s_1295;
  wire [0:0] s_1296;
  wire [0:0] s_1297;
  wire [1:0] s_1298;
  wire [3:0] s_1299;
  wire [0:0] s_1300;
  wire [0:0] s_1301;
  wire [0:0] s_1302;
  wire [0:0] s_1303;
  wire [0:0] s_1304;
  wire [0:0] s_1305;
  wire [0:0] s_1306;
  wire [1:0] s_1307;
  wire [0:0] s_1308;
  wire [0:0] s_1309;
  wire [0:0] s_1310;
  wire [1:0] s_1311;
  wire [0:0] s_1312;
  wire [0:0] s_1313;
  wire [0:0] s_1314;
  wire [0:0] s_1315;
  wire [0:0] s_1316;
  wire [0:0] s_1317;
  wire [1:0] s_1318;
  wire [0:0] s_1319;
  wire [0:0] s_1320;
  wire [0:0] s_1321;
  wire [0:0] s_1322;
  wire [0:0] s_1323;
  wire [2:0] s_1324;
  wire [0:0] s_1325;
  wire [0:0] s_1326;
  wire [1:0] s_1327;
  wire [1:0] s_1328;
  wire [1:0] s_1329;
  wire [3:0] s_1330;
  wire [0:0] s_1331;
  wire [0:0] s_1332;
  wire [2:0] s_1333;
  wire [2:0] s_1334;
  wire [2:0] s_1335;
  wire [4:0] s_1336;
  wire [0:0] s_1337;
  wire [0:0] s_1338;
  wire [3:0] s_1339;
  wire [3:0] s_1340;
  wire [3:0] s_1341;
  wire [0:0] s_1342;
  wire [5:0] s_1343;
  wire [0:0] s_1344;
  wire [0:0] s_1345;
  wire [4:0] s_1346;
  wire [0:0] s_1347;
  wire [0:0] s_1348;
  wire [3:0] s_1349;
  wire [0:0] s_1350;
  wire [0:0] s_1351;
  wire [2:0] s_1352;
  wire [0:0] s_1353;
  wire [0:0] s_1354;
  wire [1:0] s_1355;
  wire [0:0] s_1356;
  wire [0:0] s_1357;
  wire [0:0] s_1358;
  wire [1:0] s_1359;
  wire [3:0] s_1360;
  wire [7:0] s_1361;
  wire [15:0] s_1362;
  wire [31:0] s_1363;
  wire [0:0] s_1364;
  wire [0:0] s_1365;
  wire [0:0] s_1366;
  wire [0:0] s_1367;
  wire [0:0] s_1368;
  wire [0:0] s_1369;
  wire [0:0] s_1370;
  wire [1:0] s_1371;
  wire [0:0] s_1372;
  wire [0:0] s_1373;
  wire [0:0] s_1374;
  wire [1:0] s_1375;
  wire [0:0] s_1376;
  wire [0:0] s_1377;
  wire [0:0] s_1378;
  wire [0:0] s_1379;
  wire [0:0] s_1380;
  wire [0:0] s_1381;
  wire [1:0] s_1382;
  wire [0:0] s_1383;
  wire [0:0] s_1384;
  wire [0:0] s_1385;
  wire [0:0] s_1386;
  wire [0:0] s_1387;
  wire [0:0] s_1388;
  wire [2:0] s_1389;
  wire [0:0] s_1390;
  wire [0:0] s_1391;
  wire [1:0] s_1392;
  wire [0:0] s_1393;
  wire [0:0] s_1394;
  wire [0:0] s_1395;
  wire [1:0] s_1396;
  wire [3:0] s_1397;
  wire [0:0] s_1398;
  wire [0:0] s_1399;
  wire [0:0] s_1400;
  wire [0:0] s_1401;
  wire [0:0] s_1402;
  wire [0:0] s_1403;
  wire [0:0] s_1404;
  wire [1:0] s_1405;
  wire [0:0] s_1406;
  wire [0:0] s_1407;
  wire [0:0] s_1408;
  wire [1:0] s_1409;
  wire [0:0] s_1410;
  wire [0:0] s_1411;
  wire [0:0] s_1412;
  wire [0:0] s_1413;
  wire [0:0] s_1414;
  wire [0:0] s_1415;
  wire [1:0] s_1416;
  wire [0:0] s_1417;
  wire [0:0] s_1418;
  wire [0:0] s_1419;
  wire [0:0] s_1420;
  wire [0:0] s_1421;
  wire [2:0] s_1422;
  wire [0:0] s_1423;
  wire [0:0] s_1424;
  wire [1:0] s_1425;
  wire [1:0] s_1426;
  wire [1:0] s_1427;
  wire [0:0] s_1428;
  wire [3:0] s_1429;
  wire [0:0] s_1430;
  wire [0:0] s_1431;
  wire [2:0] s_1432;
  wire [0:0] s_1433;
  wire [0:0] s_1434;
  wire [1:0] s_1435;
  wire [0:0] s_1436;
  wire [0:0] s_1437;
  wire [0:0] s_1438;
  wire [1:0] s_1439;
  wire [3:0] s_1440;
  wire [7:0] s_1441;
  wire [0:0] s_1442;
  wire [0:0] s_1443;
  wire [0:0] s_1444;
  wire [0:0] s_1445;
  wire [0:0] s_1446;
  wire [0:0] s_1447;
  wire [0:0] s_1448;
  wire [1:0] s_1449;
  wire [0:0] s_1450;
  wire [0:0] s_1451;
  wire [0:0] s_1452;
  wire [1:0] s_1453;
  wire [0:0] s_1454;
  wire [0:0] s_1455;
  wire [0:0] s_1456;
  wire [0:0] s_1457;
  wire [0:0] s_1458;
  wire [0:0] s_1459;
  wire [1:0] s_1460;
  wire [0:0] s_1461;
  wire [0:0] s_1462;
  wire [0:0] s_1463;
  wire [0:0] s_1464;
  wire [0:0] s_1465;
  wire [0:0] s_1466;
  wire [2:0] s_1467;
  wire [0:0] s_1468;
  wire [0:0] s_1469;
  wire [1:0] s_1470;
  wire [0:0] s_1471;
  wire [0:0] s_1472;
  wire [0:0] s_1473;
  wire [1:0] s_1474;
  wire [3:0] s_1475;
  wire [0:0] s_1476;
  wire [0:0] s_1477;
  wire [0:0] s_1478;
  wire [0:0] s_1479;
  wire [0:0] s_1480;
  wire [0:0] s_1481;
  wire [0:0] s_1482;
  wire [1:0] s_1483;
  wire [0:0] s_1484;
  wire [0:0] s_1485;
  wire [0:0] s_1486;
  wire [1:0] s_1487;
  wire [0:0] s_1488;
  wire [0:0] s_1489;
  wire [0:0] s_1490;
  wire [0:0] s_1491;
  wire [0:0] s_1492;
  wire [0:0] s_1493;
  wire [1:0] s_1494;
  wire [0:0] s_1495;
  wire [0:0] s_1496;
  wire [0:0] s_1497;
  wire [0:0] s_1498;
  wire [0:0] s_1499;
  wire [2:0] s_1500;
  wire [0:0] s_1501;
  wire [0:0] s_1502;
  wire [1:0] s_1503;
  wire [1:0] s_1504;
  wire [1:0] s_1505;
  wire [3:0] s_1506;
  wire [0:0] s_1507;
  wire [0:0] s_1508;
  wire [2:0] s_1509;
  wire [2:0] s_1510;
  wire [2:0] s_1511;
  wire [0:0] s_1512;
  wire [4:0] s_1513;
  wire [0:0] s_1514;
  wire [0:0] s_1515;
  wire [3:0] s_1516;
  wire [0:0] s_1517;
  wire [0:0] s_1518;
  wire [2:0] s_1519;
  wire [0:0] s_1520;
  wire [0:0] s_1521;
  wire [1:0] s_1522;
  wire [0:0] s_1523;
  wire [0:0] s_1524;
  wire [0:0] s_1525;
  wire [1:0] s_1526;
  wire [3:0] s_1527;
  wire [7:0] s_1528;
  wire [15:0] s_1529;
  wire [0:0] s_1530;
  wire [0:0] s_1531;
  wire [0:0] s_1532;
  wire [0:0] s_1533;
  wire [0:0] s_1534;
  wire [0:0] s_1535;
  wire [0:0] s_1536;
  wire [1:0] s_1537;
  wire [0:0] s_1538;
  wire [0:0] s_1539;
  wire [0:0] s_1540;
  wire [1:0] s_1541;
  wire [0:0] s_1542;
  wire [0:0] s_1543;
  wire [0:0] s_1544;
  wire [0:0] s_1545;
  wire [0:0] s_1546;
  wire [0:0] s_1547;
  wire [1:0] s_1548;
  wire [0:0] s_1549;
  wire [0:0] s_1550;
  wire [0:0] s_1551;
  wire [0:0] s_1552;
  wire [0:0] s_1553;
  wire [0:0] s_1554;
  wire [2:0] s_1555;
  wire [0:0] s_1556;
  wire [0:0] s_1557;
  wire [1:0] s_1558;
  wire [0:0] s_1559;
  wire [0:0] s_1560;
  wire [0:0] s_1561;
  wire [1:0] s_1562;
  wire [3:0] s_1563;
  wire [0:0] s_1564;
  wire [0:0] s_1565;
  wire [0:0] s_1566;
  wire [0:0] s_1567;
  wire [0:0] s_1568;
  wire [0:0] s_1569;
  wire [0:0] s_1570;
  wire [1:0] s_1571;
  wire [0:0] s_1572;
  wire [0:0] s_1573;
  wire [0:0] s_1574;
  wire [1:0] s_1575;
  wire [0:0] s_1576;
  wire [0:0] s_1577;
  wire [0:0] s_1578;
  wire [0:0] s_1579;
  wire [0:0] s_1580;
  wire [0:0] s_1581;
  wire [1:0] s_1582;
  wire [0:0] s_1583;
  wire [0:0] s_1584;
  wire [0:0] s_1585;
  wire [0:0] s_1586;
  wire [0:0] s_1587;
  wire [2:0] s_1588;
  wire [0:0] s_1589;
  wire [0:0] s_1590;
  wire [1:0] s_1591;
  wire [1:0] s_1592;
  wire [1:0] s_1593;
  wire [0:0] s_1594;
  wire [3:0] s_1595;
  wire [0:0] s_1596;
  wire [0:0] s_1597;
  wire [2:0] s_1598;
  wire [0:0] s_1599;
  wire [0:0] s_1600;
  wire [1:0] s_1601;
  wire [0:0] s_1602;
  wire [0:0] s_1603;
  wire [0:0] s_1604;
  wire [1:0] s_1605;
  wire [3:0] s_1606;
  wire [7:0] s_1607;
  wire [0:0] s_1608;
  wire [0:0] s_1609;
  wire [0:0] s_1610;
  wire [0:0] s_1611;
  wire [0:0] s_1612;
  wire [0:0] s_1613;
  wire [0:0] s_1614;
  wire [1:0] s_1615;
  wire [0:0] s_1616;
  wire [0:0] s_1617;
  wire [0:0] s_1618;
  wire [1:0] s_1619;
  wire [0:0] s_1620;
  wire [0:0] s_1621;
  wire [0:0] s_1622;
  wire [0:0] s_1623;
  wire [0:0] s_1624;
  wire [0:0] s_1625;
  wire [1:0] s_1626;
  wire [0:0] s_1627;
  wire [0:0] s_1628;
  wire [0:0] s_1629;
  wire [0:0] s_1630;
  wire [0:0] s_1631;
  wire [0:0] s_1632;
  wire [2:0] s_1633;
  wire [0:0] s_1634;
  wire [0:0] s_1635;
  wire [1:0] s_1636;
  wire [0:0] s_1637;
  wire [0:0] s_1638;
  wire [0:0] s_1639;
  wire [1:0] s_1640;
  wire [3:0] s_1641;
  wire [0:0] s_1642;
  wire [0:0] s_1643;
  wire [0:0] s_1644;
  wire [0:0] s_1645;
  wire [0:0] s_1646;
  wire [0:0] s_1647;
  wire [0:0] s_1648;
  wire [1:0] s_1649;
  wire [0:0] s_1650;
  wire [0:0] s_1651;
  wire [0:0] s_1652;
  wire [1:0] s_1653;
  wire [0:0] s_1654;
  wire [0:0] s_1655;
  wire [0:0] s_1656;
  wire [0:0] s_1657;
  wire [0:0] s_1658;
  wire [0:0] s_1659;
  wire [1:0] s_1660;
  wire [0:0] s_1661;
  wire [0:0] s_1662;
  wire [0:0] s_1663;
  wire [0:0] s_1664;
  wire [0:0] s_1665;
  wire [2:0] s_1666;
  wire [0:0] s_1667;
  wire [0:0] s_1668;
  wire [1:0] s_1669;
  wire [1:0] s_1670;
  wire [1:0] s_1671;
  wire [3:0] s_1672;
  wire [0:0] s_1673;
  wire [0:0] s_1674;
  wire [2:0] s_1675;
  wire [2:0] s_1676;
  wire [2:0] s_1677;
  wire [4:0] s_1678;
  wire [0:0] s_1679;
  wire [0:0] s_1680;
  wire [3:0] s_1681;
  wire [3:0] s_1682;
  wire [3:0] s_1683;
  wire [5:0] s_1684;
  wire [0:0] s_1685;
  wire [0:0] s_1686;
  wire [4:0] s_1687;
  wire [4:0] s_1688;
  wire [4:0] s_1689;
  wire [12:0] s_1690;
  wire [12:0] s_1691;
  wire [12:0] s_1692;
  wire [10:0] s_1693;
  wire [10:0] s_1694;
  wire [12:0] s_1695;
  wire [0:0] s_1696;
  wire [12:0] s_1697;
  wire [12:0] s_1698;
  wire [1:0] s_1699;
  wire [0:0] s_1700;
  wire [55:0] s_1701;
  wire [0:0] s_1702;
  wire [0:0] s_1703;
  wire [56:0] s_1704;
  wire [56:0] s_1705;
  wire [56:0] s_1706;
  wire [56:0] s_1707;
  wire [56:0] s_1708;
  wire [56:0] s_1709;
  wire [0:0] s_1710;
  wire [0:0] s_1711;
  wire [55:0] s_1712;
  wire [0:0] s_1713;
  wire [55:0] s_1714;
  wire [0:0] s_1715;
  wire [0:0] s_1716;
  wire [56:0] s_1717;
  wire [56:0] s_1718;
  wire [56:0] s_1719;
  wire [56:0] s_1720;
  wire [56:0] s_1721;
  wire [56:0] s_1722;
  wire [0:0] s_1723;
  wire [0:0] s_1724;
  wire [55:0] s_1725;
  wire [0:0] s_1726;
  wire [55:0] s_1727;
  wire [0:0] s_1728;
  wire [0:0] s_1729;
  wire [56:0] s_1730;
  wire [56:0] s_1731;
  wire [56:0] s_1732;
  wire [56:0] s_1733;
  wire [56:0] s_1734;
  wire [56:0] s_1735;
  wire [0:0] s_1736;
  wire [0:0] s_1737;
  wire [55:0] s_1738;
  wire [0:0] s_1739;
  wire [55:0] s_1740;
  wire [0:0] s_1741;
  wire [0:0] s_1742;
  wire [56:0] s_1743;
  wire [56:0] s_1744;
  wire [56:0] s_1745;
  wire [56:0] s_1746;
  wire [56:0] s_1747;
  wire [56:0] s_1748;
  wire [0:0] s_1749;
  wire [0:0] s_1750;
  wire [55:0] s_1751;
  wire [0:0] s_1752;
  wire [55:0] s_1753;
  wire [0:0] s_1754;
  wire [0:0] s_1755;
  wire [56:0] s_1756;
  wire [56:0] s_1757;
  wire [56:0] s_1758;
  wire [56:0] s_1759;
  wire [56:0] s_1760;
  wire [56:0] s_1761;
  wire [0:0] s_1762;
  wire [0:0] s_1763;
  wire [55:0] s_1764;
  wire [0:0] s_1765;
  wire [55:0] s_1766;
  wire [0:0] s_1767;
  wire [0:0] s_1768;
  wire [56:0] s_1769;
  wire [56:0] s_1770;
  wire [56:0] s_1771;
  wire [56:0] s_1772;
  wire [56:0] s_1773;
  wire [56:0] s_1774;
  wire [0:0] s_1775;
  wire [0:0] s_1776;
  wire [55:0] s_1777;
  wire [0:0] s_1778;
  wire [55:0] s_1779;
  wire [0:0] s_1780;
  wire [0:0] s_1781;
  wire [56:0] s_1782;
  wire [56:0] s_1783;
  wire [56:0] s_1784;
  wire [56:0] s_1785;
  wire [56:0] s_1786;
  wire [56:0] s_1787;
  wire [0:0] s_1788;
  wire [0:0] s_1789;
  wire [55:0] s_1790;
  wire [0:0] s_1791;
  wire [55:0] s_1792;
  wire [0:0] s_1793;
  wire [0:0] s_1794;
  wire [56:0] s_1795;
  wire [56:0] s_1796;
  wire [56:0] s_1797;
  wire [56:0] s_1798;
  wire [56:0] s_1799;
  wire [56:0] s_1800;
  wire [0:0] s_1801;
  wire [0:0] s_1802;
  wire [55:0] s_1803;
  wire [0:0] s_1804;
  wire [55:0] s_1805;
  wire [0:0] s_1806;
  wire [0:0] s_1807;
  wire [56:0] s_1808;
  wire [56:0] s_1809;
  wire [56:0] s_1810;
  wire [56:0] s_1811;
  wire [56:0] s_1812;
  wire [56:0] s_1813;
  wire [0:0] s_1814;
  wire [0:0] s_1815;
  wire [55:0] s_1816;
  wire [0:0] s_1817;
  wire [55:0] s_1818;
  wire [0:0] s_1819;
  wire [0:0] s_1820;
  wire [56:0] s_1821;
  wire [56:0] s_1822;
  wire [56:0] s_1823;
  wire [56:0] s_1824;
  wire [56:0] s_1825;
  wire [56:0] s_1826;
  wire [0:0] s_1827;
  wire [0:0] s_1828;
  wire [55:0] s_1829;
  wire [0:0] s_1830;
  wire [55:0] s_1831;
  wire [0:0] s_1832;
  wire [0:0] s_1833;
  wire [56:0] s_1834;
  wire [56:0] s_1835;
  wire [56:0] s_1836;
  wire [56:0] s_1837;
  wire [56:0] s_1838;
  wire [56:0] s_1839;
  wire [0:0] s_1840;
  wire [0:0] s_1841;
  wire [55:0] s_1842;
  wire [0:0] s_1843;
  wire [55:0] s_1844;
  wire [0:0] s_1845;
  wire [0:0] s_1846;
  wire [56:0] s_1847;
  wire [56:0] s_1848;
  wire [56:0] s_1849;
  wire [56:0] s_1850;
  wire [56:0] s_1851;
  wire [56:0] s_1852;
  wire [0:0] s_1853;
  wire [0:0] s_1854;
  wire [55:0] s_1855;
  wire [0:0] s_1856;
  wire [55:0] s_1857;
  wire [0:0] s_1858;
  wire [0:0] s_1859;
  wire [56:0] s_1860;
  wire [56:0] s_1861;
  wire [56:0] s_1862;
  wire [56:0] s_1863;
  wire [56:0] s_1864;
  wire [56:0] s_1865;
  wire [0:0] s_1866;
  wire [0:0] s_1867;
  wire [55:0] s_1868;
  wire [0:0] s_1869;
  wire [55:0] s_1870;
  wire [0:0] s_1871;
  wire [0:0] s_1872;
  wire [56:0] s_1873;
  wire [56:0] s_1874;
  wire [56:0] s_1875;
  wire [56:0] s_1876;
  wire [56:0] s_1877;
  wire [56:0] s_1878;
  wire [0:0] s_1879;
  wire [0:0] s_1880;
  wire [55:0] s_1881;
  wire [0:0] s_1882;
  wire [55:0] s_1883;
  wire [0:0] s_1884;
  wire [0:0] s_1885;
  wire [56:0] s_1886;
  wire [56:0] s_1887;
  wire [56:0] s_1888;
  wire [56:0] s_1889;
  wire [56:0] s_1890;
  wire [56:0] s_1891;
  wire [0:0] s_1892;
  wire [0:0] s_1893;
  wire [55:0] s_1894;
  wire [0:0] s_1895;
  wire [55:0] s_1896;
  wire [0:0] s_1897;
  wire [0:0] s_1898;
  wire [56:0] s_1899;
  wire [56:0] s_1900;
  wire [56:0] s_1901;
  wire [56:0] s_1902;
  wire [56:0] s_1903;
  wire [56:0] s_1904;
  wire [0:0] s_1905;
  wire [0:0] s_1906;
  wire [55:0] s_1907;
  wire [0:0] s_1908;
  wire [55:0] s_1909;
  wire [0:0] s_1910;
  wire [0:0] s_1911;
  wire [56:0] s_1912;
  wire [56:0] s_1913;
  wire [56:0] s_1914;
  wire [56:0] s_1915;
  wire [56:0] s_1916;
  wire [56:0] s_1917;
  wire [0:0] s_1918;
  wire [0:0] s_1919;
  wire [55:0] s_1920;
  wire [0:0] s_1921;
  wire [55:0] s_1922;
  wire [0:0] s_1923;
  wire [0:0] s_1924;
  wire [56:0] s_1925;
  wire [56:0] s_1926;
  wire [56:0] s_1927;
  wire [56:0] s_1928;
  wire [56:0] s_1929;
  wire [56:0] s_1930;
  wire [0:0] s_1931;
  wire [0:0] s_1932;
  wire [55:0] s_1933;
  wire [0:0] s_1934;
  wire [55:0] s_1935;
  wire [0:0] s_1936;
  wire [0:0] s_1937;
  wire [56:0] s_1938;
  wire [56:0] s_1939;
  wire [56:0] s_1940;
  wire [56:0] s_1941;
  wire [56:0] s_1942;
  wire [56:0] s_1943;
  wire [0:0] s_1944;
  wire [0:0] s_1945;
  wire [55:0] s_1946;
  wire [0:0] s_1947;
  wire [55:0] s_1948;
  wire [0:0] s_1949;
  wire [0:0] s_1950;
  wire [56:0] s_1951;
  wire [56:0] s_1952;
  wire [56:0] s_1953;
  wire [56:0] s_1954;
  wire [56:0] s_1955;
  wire [56:0] s_1956;
  wire [0:0] s_1957;
  wire [0:0] s_1958;
  wire [55:0] s_1959;
  wire [0:0] s_1960;
  wire [55:0] s_1961;
  wire [0:0] s_1962;
  wire [0:0] s_1963;
  wire [56:0] s_1964;
  wire [56:0] s_1965;
  wire [56:0] s_1966;
  wire [56:0] s_1967;
  wire [56:0] s_1968;
  wire [56:0] s_1969;
  wire [0:0] s_1970;
  wire [0:0] s_1971;
  wire [55:0] s_1972;
  wire [0:0] s_1973;
  wire [55:0] s_1974;
  wire [0:0] s_1975;
  wire [0:0] s_1976;
  wire [56:0] s_1977;
  wire [56:0] s_1978;
  wire [56:0] s_1979;
  wire [56:0] s_1980;
  wire [56:0] s_1981;
  wire [56:0] s_1982;
  wire [0:0] s_1983;
  wire [0:0] s_1984;
  wire [55:0] s_1985;
  wire [0:0] s_1986;
  wire [55:0] s_1987;
  wire [0:0] s_1988;
  wire [0:0] s_1989;
  wire [56:0] s_1990;
  wire [56:0] s_1991;
  wire [56:0] s_1992;
  wire [56:0] s_1993;
  wire [56:0] s_1994;
  wire [56:0] s_1995;
  wire [0:0] s_1996;
  wire [0:0] s_1997;
  wire [55:0] s_1998;
  wire [0:0] s_1999;
  wire [55:0] s_2000;
  wire [0:0] s_2001;
  wire [0:0] s_2002;
  wire [56:0] s_2003;
  wire [56:0] s_2004;
  wire [56:0] s_2005;
  wire [56:0] s_2006;
  wire [56:0] s_2007;
  wire [56:0] s_2008;
  wire [0:0] s_2009;
  wire [0:0] s_2010;
  wire [55:0] s_2011;
  wire [0:0] s_2012;
  wire [55:0] s_2013;
  wire [0:0] s_2014;
  wire [0:0] s_2015;
  wire [56:0] s_2016;
  wire [56:0] s_2017;
  wire [56:0] s_2018;
  wire [56:0] s_2019;
  wire [56:0] s_2020;
  wire [56:0] s_2021;
  wire [0:0] s_2022;
  wire [0:0] s_2023;
  wire [55:0] s_2024;
  wire [0:0] s_2025;
  wire [55:0] s_2026;
  wire [0:0] s_2027;
  wire [0:0] s_2028;
  wire [56:0] s_2029;
  wire [56:0] s_2030;
  wire [56:0] s_2031;
  wire [56:0] s_2032;
  wire [56:0] s_2033;
  wire [56:0] s_2034;
  wire [0:0] s_2035;
  wire [0:0] s_2036;
  wire [55:0] s_2037;
  wire [0:0] s_2038;
  wire [55:0] s_2039;
  wire [0:0] s_2040;
  wire [0:0] s_2041;
  wire [56:0] s_2042;
  wire [56:0] s_2043;
  wire [56:0] s_2044;
  wire [56:0] s_2045;
  wire [56:0] s_2046;
  wire [56:0] s_2047;
  wire [0:0] s_2048;
  wire [0:0] s_2049;
  wire [55:0] s_2050;
  wire [0:0] s_2051;
  wire [55:0] s_2052;
  wire [0:0] s_2053;
  wire [0:0] s_2054;
  wire [56:0] s_2055;
  wire [56:0] s_2056;
  wire [56:0] s_2057;
  wire [56:0] s_2058;
  wire [56:0] s_2059;
  wire [56:0] s_2060;
  wire [0:0] s_2061;
  wire [0:0] s_2062;
  wire [55:0] s_2063;
  wire [0:0] s_2064;
  wire [55:0] s_2065;
  wire [0:0] s_2066;
  wire [0:0] s_2067;
  wire [56:0] s_2068;
  wire [56:0] s_2069;
  wire [56:0] s_2070;
  wire [56:0] s_2071;
  wire [56:0] s_2072;
  wire [56:0] s_2073;
  wire [0:0] s_2074;
  wire [0:0] s_2075;
  wire [55:0] s_2076;
  wire [0:0] s_2077;
  wire [55:0] s_2078;
  wire [0:0] s_2079;
  wire [0:0] s_2080;
  wire [56:0] s_2081;
  wire [56:0] s_2082;
  wire [56:0] s_2083;
  wire [56:0] s_2084;
  wire [56:0] s_2085;
  wire [56:0] s_2086;
  wire [0:0] s_2087;
  wire [0:0] s_2088;
  wire [55:0] s_2089;
  wire [0:0] s_2090;
  wire [55:0] s_2091;
  wire [0:0] s_2092;
  wire [0:0] s_2093;
  wire [56:0] s_2094;
  wire [56:0] s_2095;
  wire [56:0] s_2096;
  wire [56:0] s_2097;
  wire [56:0] s_2098;
  wire [56:0] s_2099;
  wire [0:0] s_2100;
  wire [0:0] s_2101;
  wire [55:0] s_2102;
  wire [0:0] s_2103;
  wire [55:0] s_2104;
  wire [0:0] s_2105;
  wire [0:0] s_2106;
  wire [56:0] s_2107;
  wire [56:0] s_2108;
  wire [56:0] s_2109;
  wire [56:0] s_2110;
  wire [56:0] s_2111;
  wire [56:0] s_2112;
  wire [0:0] s_2113;
  wire [0:0] s_2114;
  wire [55:0] s_2115;
  wire [0:0] s_2116;
  wire [55:0] s_2117;
  wire [0:0] s_2118;
  wire [0:0] s_2119;
  wire [56:0] s_2120;
  wire [56:0] s_2121;
  wire [56:0] s_2122;
  wire [56:0] s_2123;
  wire [56:0] s_2124;
  wire [56:0] s_2125;
  wire [0:0] s_2126;
  wire [0:0] s_2127;
  wire [55:0] s_2128;
  wire [0:0] s_2129;
  wire [55:0] s_2130;
  wire [0:0] s_2131;
  wire [0:0] s_2132;
  wire [56:0] s_2133;
  wire [56:0] s_2134;
  wire [56:0] s_2135;
  wire [56:0] s_2136;
  wire [56:0] s_2137;
  wire [56:0] s_2138;
  wire [0:0] s_2139;
  wire [0:0] s_2140;
  wire [55:0] s_2141;
  wire [0:0] s_2142;
  wire [55:0] s_2143;
  wire [0:0] s_2144;
  wire [0:0] s_2145;
  wire [56:0] s_2146;
  wire [56:0] s_2147;
  wire [56:0] s_2148;
  wire [56:0] s_2149;
  wire [56:0] s_2150;
  wire [56:0] s_2151;
  wire [0:0] s_2152;
  wire [0:0] s_2153;
  wire [55:0] s_2154;
  wire [0:0] s_2155;
  wire [55:0] s_2156;
  wire [0:0] s_2157;
  wire [0:0] s_2158;
  wire [56:0] s_2159;
  wire [56:0] s_2160;
  wire [56:0] s_2161;
  wire [56:0] s_2162;
  wire [56:0] s_2163;
  wire [56:0] s_2164;
  wire [0:0] s_2165;
  wire [0:0] s_2166;
  wire [55:0] s_2167;
  wire [0:0] s_2168;
  wire [55:0] s_2169;
  wire [0:0] s_2170;
  wire [0:0] s_2171;
  wire [56:0] s_2172;
  wire [56:0] s_2173;
  wire [56:0] s_2174;
  wire [56:0] s_2175;
  wire [56:0] s_2176;
  wire [56:0] s_2177;
  wire [0:0] s_2178;
  wire [0:0] s_2179;
  wire [55:0] s_2180;
  wire [0:0] s_2181;
  wire [55:0] s_2182;
  wire [0:0] s_2183;
  wire [0:0] s_2184;
  wire [56:0] s_2185;
  wire [56:0] s_2186;
  wire [56:0] s_2187;
  wire [56:0] s_2188;
  wire [56:0] s_2189;
  wire [56:0] s_2190;
  wire [0:0] s_2191;
  wire [0:0] s_2192;
  wire [55:0] s_2193;
  wire [0:0] s_2194;
  wire [55:0] s_2195;
  wire [0:0] s_2196;
  wire [0:0] s_2197;
  wire [56:0] s_2198;
  wire [56:0] s_2199;
  wire [56:0] s_2200;
  wire [56:0] s_2201;
  wire [56:0] s_2202;
  wire [56:0] s_2203;
  wire [0:0] s_2204;
  wire [0:0] s_2205;
  wire [55:0] s_2206;
  wire [0:0] s_2207;
  wire [55:0] s_2208;
  wire [0:0] s_2209;
  wire [0:0] s_2210;
  wire [56:0] s_2211;
  wire [56:0] s_2212;
  wire [56:0] s_2213;
  wire [56:0] s_2214;
  wire [56:0] s_2215;
  wire [56:0] s_2216;
  wire [0:0] s_2217;
  wire [0:0] s_2218;
  wire [55:0] s_2219;
  wire [0:0] s_2220;
  wire [55:0] s_2221;
  wire [0:0] s_2222;
  wire [0:0] s_2223;
  wire [56:0] s_2224;
  wire [56:0] s_2225;
  wire [56:0] s_2226;
  wire [56:0] s_2227;
  wire [56:0] s_2228;
  wire [56:0] s_2229;
  wire [0:0] s_2230;
  wire [0:0] s_2231;
  wire [55:0] s_2232;
  wire [0:0] s_2233;
  wire [55:0] s_2234;
  wire [0:0] s_2235;
  wire [0:0] s_2236;
  wire [56:0] s_2237;
  wire [56:0] s_2238;
  wire [56:0] s_2239;
  wire [56:0] s_2240;
  wire [56:0] s_2241;
  wire [56:0] s_2242;
  wire [0:0] s_2243;
  wire [0:0] s_2244;
  wire [55:0] s_2245;
  wire [0:0] s_2246;
  wire [55:0] s_2247;
  wire [0:0] s_2248;
  wire [0:0] s_2249;
  wire [56:0] s_2250;
  wire [56:0] s_2251;
  wire [56:0] s_2252;
  wire [56:0] s_2253;
  wire [56:0] s_2254;
  wire [56:0] s_2255;
  wire [0:0] s_2256;
  wire [0:0] s_2257;
  wire [55:0] s_2258;
  wire [0:0] s_2259;
  wire [55:0] s_2260;
  wire [0:0] s_2261;
  wire [0:0] s_2262;
  wire [56:0] s_2263;
  wire [56:0] s_2264;
  wire [56:0] s_2265;
  wire [56:0] s_2266;
  wire [56:0] s_2267;
  wire [56:0] s_2268;
  wire [0:0] s_2269;
  wire [0:0] s_2270;
  wire [55:0] s_2271;
  wire [0:0] s_2272;
  wire [55:0] s_2273;
  wire [0:0] s_2274;
  wire [0:0] s_2275;
  wire [56:0] s_2276;
  wire [56:0] s_2277;
  wire [56:0] s_2278;
  wire [56:0] s_2279;
  wire [56:0] s_2280;
  wire [56:0] s_2281;
  wire [0:0] s_2282;
  wire [0:0] s_2283;
  wire [55:0] s_2284;
  wire [0:0] s_2285;
  wire [55:0] s_2286;
  wire [0:0] s_2287;
  wire [0:0] s_2288;
  wire [56:0] s_2289;
  wire [56:0] s_2290;
  wire [56:0] s_2291;
  wire [56:0] s_2292;
  wire [56:0] s_2293;
  wire [56:0] s_2294;
  wire [0:0] s_2295;
  wire [0:0] s_2296;
  wire [55:0] s_2297;
  wire [0:0] s_2298;
  wire [55:0] s_2299;
  wire [0:0] s_2300;
  wire [0:0] s_2301;
  wire [56:0] s_2302;
  wire [56:0] s_2303;
  wire [56:0] s_2304;
  wire [56:0] s_2305;
  wire [56:0] s_2306;
  wire [56:0] s_2307;
  wire [0:0] s_2308;
  wire [0:0] s_2309;
  wire [55:0] s_2310;
  wire [0:0] s_2311;
  wire [55:0] s_2312;
  wire [0:0] s_2313;
  wire [0:0] s_2314;
  wire [56:0] s_2315;
  wire [56:0] s_2316;
  wire [56:0] s_2317;
  wire [56:0] s_2318;
  wire [56:0] s_2319;
  wire [56:0] s_2320;
  wire [0:0] s_2321;
  wire [0:0] s_2322;
  wire [55:0] s_2323;
  wire [0:0] s_2324;
  wire [55:0] s_2325;
  wire [0:0] s_2326;
  wire [0:0] s_2327;
  wire [56:0] s_2328;
  wire [56:0] s_2329;
  wire [56:0] s_2330;
  wire [56:0] s_2331;
  wire [56:0] s_2332;
  wire [56:0] s_2333;
  wire [0:0] s_2334;
  wire [0:0] s_2335;
  wire [55:0] s_2336;
  wire [0:0] s_2337;
  wire [55:0] s_2338;
  wire [0:0] s_2339;
  wire [0:0] s_2340;
  wire [56:0] s_2341;
  wire [56:0] s_2342;
  wire [56:0] s_2343;
  wire [56:0] s_2344;
  wire [56:0] s_2345;
  wire [56:0] s_2346;
  wire [0:0] s_2347;
  wire [0:0] s_2348;
  wire [55:0] s_2349;
  wire [0:0] s_2350;
  wire [55:0] s_2351;
  wire [0:0] s_2352;
  wire [0:0] s_2353;
  wire [56:0] s_2354;
  wire [56:0] s_2355;
  wire [56:0] s_2356;
  wire [56:0] s_2357;
  wire [56:0] s_2358;
  wire [56:0] s_2359;
  wire [0:0] s_2360;
  wire [0:0] s_2361;
  wire [55:0] s_2362;
  wire [0:0] s_2363;
  wire [55:0] s_2364;
  wire [0:0] s_2365;
  wire [0:0] s_2366;
  wire [56:0] s_2367;
  wire [56:0] s_2368;
  wire [56:0] s_2369;
  wire [56:0] s_2370;
  wire [56:0] s_2371;
  wire [56:0] s_2372;
  wire [0:0] s_2373;
  wire [0:0] s_2374;
  wire [55:0] s_2375;
  wire [0:0] s_2376;
  wire [55:0] s_2377;
  wire [0:0] s_2378;
  wire [0:0] s_2379;
  wire [56:0] s_2380;
  wire [56:0] s_2381;
  wire [56:0] s_2382;
  wire [56:0] s_2383;
  wire [56:0] s_2384;
  wire [56:0] s_2385;
  wire [0:0] s_2386;
  wire [0:0] s_2387;
  wire [55:0] s_2388;
  wire [0:0] s_2389;
  wire [55:0] s_2390;
  wire [0:0] s_2391;
  wire [0:0] s_2392;
  wire [56:0] s_2393;
  wire [56:0] s_2394;
  wire [56:0] s_2395;
  wire [56:0] s_2396;
  wire [56:0] s_2397;
  wire [56:0] s_2398;
  wire [0:0] s_2399;
  wire [0:0] s_2400;
  wire [55:0] s_2401;
  wire [0:0] s_2402;
  wire [55:0] s_2403;
  wire [0:0] s_2404;
  wire [0:0] s_2405;
  wire [56:0] s_2406;
  wire [56:0] s_2407;
  wire [56:0] s_2408;
  wire [56:0] s_2409;
  wire [56:0] s_2410;
  wire [56:0] s_2411;
  wire [0:0] s_2412;
  wire [0:0] s_2413;
  wire [55:0] s_2414;
  wire [12:0] s_2415;
  wire [12:0] s_2416;
  wire [12:0] s_2417;
  wire [0:0] s_2418;
  wire [12:0] s_2419;
  wire [12:0] s_2420;
  wire [12:0] s_2421;
  wire [12:0] s_2422;
  wire [12:0] s_2423;
  wire [12:0] s_2424;
  wire [12:0] s_2425;
  wire [12:0] s_2426;
  wire [12:0] s_2427;
  wire [12:0] s_2428;
  wire [12:0] s_2429;
  wire [0:0] s_2430;
  wire [12:0] s_2431;
  wire [12:0] s_2432;
  wire [6:0] s_2433;
  wire [6:0] s_2434;
  wire [0:0] s_2435;
  wire [0:0] s_2436;
  wire [5:0] s_2437;
  wire [0:0] s_2438;
  wire [0:0] s_2439;
  wire [4:0] s_2440;
  wire [0:0] s_2441;
  wire [0:0] s_2442;
  wire [3:0] s_2443;
  wire [0:0] s_2444;
  wire [0:0] s_2445;
  wire [2:0] s_2446;
  wire [0:0] s_2447;
  wire [0:0] s_2448;
  wire [1:0] s_2449;
  wire [0:0] s_2450;
  wire [0:0] s_2451;
  wire [0:0] s_2452;
  wire [1:0] s_2453;
  wire [3:0] s_2454;
  wire [7:0] s_2455;
  wire [15:0] s_2456;
  wire [31:0] s_2457;
  wire [63:0] s_2458;
  wire [62:0] s_2459;
  wire [61:0] s_2460;
  wire [60:0] s_2461;
  wire [59:0] s_2462;
  wire [58:0] s_2463;
  wire [57:0] s_2464;
  wire [56:0] s_2465;
  wire [0:0] s_2466;
  wire [0:0] s_2467;
  wire [0:0] s_2468;
  wire [0:0] s_2469;
  wire [0:0] s_2470;
  wire [0:0] s_2471;
  wire [0:0] s_2472;
  wire [0:0] s_2473;
  wire [0:0] s_2474;
  wire [0:0] s_2475;
  wire [0:0] s_2476;
  wire [0:0] s_2477;
  wire [0:0] s_2478;
  wire [0:0] s_2479;
  wire [0:0] s_2480;
  wire [1:0] s_2481;
  wire [0:0] s_2482;
  wire [0:0] s_2483;
  wire [0:0] s_2484;
  wire [1:0] s_2485;
  wire [0:0] s_2486;
  wire [0:0] s_2487;
  wire [0:0] s_2488;
  wire [0:0] s_2489;
  wire [0:0] s_2490;
  wire [0:0] s_2491;
  wire [1:0] s_2492;
  wire [0:0] s_2493;
  wire [0:0] s_2494;
  wire [0:0] s_2495;
  wire [0:0] s_2496;
  wire [0:0] s_2497;
  wire [0:0] s_2498;
  wire [2:0] s_2499;
  wire [0:0] s_2500;
  wire [0:0] s_2501;
  wire [1:0] s_2502;
  wire [0:0] s_2503;
  wire [0:0] s_2504;
  wire [0:0] s_2505;
  wire [1:0] s_2506;
  wire [3:0] s_2507;
  wire [0:0] s_2508;
  wire [0:0] s_2509;
  wire [0:0] s_2510;
  wire [0:0] s_2511;
  wire [0:0] s_2512;
  wire [0:0] s_2513;
  wire [0:0] s_2514;
  wire [1:0] s_2515;
  wire [0:0] s_2516;
  wire [0:0] s_2517;
  wire [0:0] s_2518;
  wire [1:0] s_2519;
  wire [0:0] s_2520;
  wire [0:0] s_2521;
  wire [0:0] s_2522;
  wire [0:0] s_2523;
  wire [0:0] s_2524;
  wire [0:0] s_2525;
  wire [1:0] s_2526;
  wire [0:0] s_2527;
  wire [0:0] s_2528;
  wire [0:0] s_2529;
  wire [0:0] s_2530;
  wire [0:0] s_2531;
  wire [2:0] s_2532;
  wire [0:0] s_2533;
  wire [0:0] s_2534;
  wire [1:0] s_2535;
  wire [1:0] s_2536;
  wire [1:0] s_2537;
  wire [0:0] s_2538;
  wire [3:0] s_2539;
  wire [0:0] s_2540;
  wire [0:0] s_2541;
  wire [2:0] s_2542;
  wire [0:0] s_2543;
  wire [0:0] s_2544;
  wire [1:0] s_2545;
  wire [0:0] s_2546;
  wire [0:0] s_2547;
  wire [0:0] s_2548;
  wire [1:0] s_2549;
  wire [3:0] s_2550;
  wire [7:0] s_2551;
  wire [0:0] s_2552;
  wire [0:0] s_2553;
  wire [0:0] s_2554;
  wire [0:0] s_2555;
  wire [0:0] s_2556;
  wire [0:0] s_2557;
  wire [0:0] s_2558;
  wire [1:0] s_2559;
  wire [0:0] s_2560;
  wire [0:0] s_2561;
  wire [0:0] s_2562;
  wire [1:0] s_2563;
  wire [0:0] s_2564;
  wire [0:0] s_2565;
  wire [0:0] s_2566;
  wire [0:0] s_2567;
  wire [0:0] s_2568;
  wire [0:0] s_2569;
  wire [1:0] s_2570;
  wire [0:0] s_2571;
  wire [0:0] s_2572;
  wire [0:0] s_2573;
  wire [0:0] s_2574;
  wire [0:0] s_2575;
  wire [0:0] s_2576;
  wire [2:0] s_2577;
  wire [0:0] s_2578;
  wire [0:0] s_2579;
  wire [1:0] s_2580;
  wire [0:0] s_2581;
  wire [0:0] s_2582;
  wire [0:0] s_2583;
  wire [1:0] s_2584;
  wire [3:0] s_2585;
  wire [0:0] s_2586;
  wire [0:0] s_2587;
  wire [0:0] s_2588;
  wire [0:0] s_2589;
  wire [0:0] s_2590;
  wire [0:0] s_2591;
  wire [0:0] s_2592;
  wire [1:0] s_2593;
  wire [0:0] s_2594;
  wire [0:0] s_2595;
  wire [0:0] s_2596;
  wire [1:0] s_2597;
  wire [0:0] s_2598;
  wire [0:0] s_2599;
  wire [0:0] s_2600;
  wire [0:0] s_2601;
  wire [0:0] s_2602;
  wire [0:0] s_2603;
  wire [1:0] s_2604;
  wire [0:0] s_2605;
  wire [0:0] s_2606;
  wire [0:0] s_2607;
  wire [0:0] s_2608;
  wire [0:0] s_2609;
  wire [2:0] s_2610;
  wire [0:0] s_2611;
  wire [0:0] s_2612;
  wire [1:0] s_2613;
  wire [1:0] s_2614;
  wire [1:0] s_2615;
  wire [3:0] s_2616;
  wire [0:0] s_2617;
  wire [0:0] s_2618;
  wire [2:0] s_2619;
  wire [2:0] s_2620;
  wire [2:0] s_2621;
  wire [0:0] s_2622;
  wire [4:0] s_2623;
  wire [0:0] s_2624;
  wire [0:0] s_2625;
  wire [3:0] s_2626;
  wire [0:0] s_2627;
  wire [0:0] s_2628;
  wire [2:0] s_2629;
  wire [0:0] s_2630;
  wire [0:0] s_2631;
  wire [1:0] s_2632;
  wire [0:0] s_2633;
  wire [0:0] s_2634;
  wire [0:0] s_2635;
  wire [1:0] s_2636;
  wire [3:0] s_2637;
  wire [7:0] s_2638;
  wire [15:0] s_2639;
  wire [0:0] s_2640;
  wire [0:0] s_2641;
  wire [0:0] s_2642;
  wire [0:0] s_2643;
  wire [0:0] s_2644;
  wire [0:0] s_2645;
  wire [0:0] s_2646;
  wire [1:0] s_2647;
  wire [0:0] s_2648;
  wire [0:0] s_2649;
  wire [0:0] s_2650;
  wire [1:0] s_2651;
  wire [0:0] s_2652;
  wire [0:0] s_2653;
  wire [0:0] s_2654;
  wire [0:0] s_2655;
  wire [0:0] s_2656;
  wire [0:0] s_2657;
  wire [1:0] s_2658;
  wire [0:0] s_2659;
  wire [0:0] s_2660;
  wire [0:0] s_2661;
  wire [0:0] s_2662;
  wire [0:0] s_2663;
  wire [0:0] s_2664;
  wire [2:0] s_2665;
  wire [0:0] s_2666;
  wire [0:0] s_2667;
  wire [1:0] s_2668;
  wire [0:0] s_2669;
  wire [0:0] s_2670;
  wire [0:0] s_2671;
  wire [1:0] s_2672;
  wire [3:0] s_2673;
  wire [0:0] s_2674;
  wire [0:0] s_2675;
  wire [0:0] s_2676;
  wire [0:0] s_2677;
  wire [0:0] s_2678;
  wire [0:0] s_2679;
  wire [0:0] s_2680;
  wire [1:0] s_2681;
  wire [0:0] s_2682;
  wire [0:0] s_2683;
  wire [0:0] s_2684;
  wire [1:0] s_2685;
  wire [0:0] s_2686;
  wire [0:0] s_2687;
  wire [0:0] s_2688;
  wire [0:0] s_2689;
  wire [0:0] s_2690;
  wire [0:0] s_2691;
  wire [1:0] s_2692;
  wire [0:0] s_2693;
  wire [0:0] s_2694;
  wire [0:0] s_2695;
  wire [0:0] s_2696;
  wire [0:0] s_2697;
  wire [2:0] s_2698;
  wire [0:0] s_2699;
  wire [0:0] s_2700;
  wire [1:0] s_2701;
  wire [1:0] s_2702;
  wire [1:0] s_2703;
  wire [0:0] s_2704;
  wire [3:0] s_2705;
  wire [0:0] s_2706;
  wire [0:0] s_2707;
  wire [2:0] s_2708;
  wire [0:0] s_2709;
  wire [0:0] s_2710;
  wire [1:0] s_2711;
  wire [0:0] s_2712;
  wire [0:0] s_2713;
  wire [0:0] s_2714;
  wire [1:0] s_2715;
  wire [3:0] s_2716;
  wire [7:0] s_2717;
  wire [0:0] s_2718;
  wire [0:0] s_2719;
  wire [0:0] s_2720;
  wire [0:0] s_2721;
  wire [0:0] s_2722;
  wire [0:0] s_2723;
  wire [0:0] s_2724;
  wire [1:0] s_2725;
  wire [0:0] s_2726;
  wire [0:0] s_2727;
  wire [0:0] s_2728;
  wire [1:0] s_2729;
  wire [0:0] s_2730;
  wire [0:0] s_2731;
  wire [0:0] s_2732;
  wire [0:0] s_2733;
  wire [0:0] s_2734;
  wire [0:0] s_2735;
  wire [1:0] s_2736;
  wire [0:0] s_2737;
  wire [0:0] s_2738;
  wire [0:0] s_2739;
  wire [0:0] s_2740;
  wire [0:0] s_2741;
  wire [0:0] s_2742;
  wire [2:0] s_2743;
  wire [0:0] s_2744;
  wire [0:0] s_2745;
  wire [1:0] s_2746;
  wire [0:0] s_2747;
  wire [0:0] s_2748;
  wire [0:0] s_2749;
  wire [1:0] s_2750;
  wire [3:0] s_2751;
  wire [0:0] s_2752;
  wire [0:0] s_2753;
  wire [0:0] s_2754;
  wire [0:0] s_2755;
  wire [0:0] s_2756;
  wire [0:0] s_2757;
  wire [0:0] s_2758;
  wire [1:0] s_2759;
  wire [0:0] s_2760;
  wire [0:0] s_2761;
  wire [0:0] s_2762;
  wire [1:0] s_2763;
  wire [0:0] s_2764;
  wire [0:0] s_2765;
  wire [0:0] s_2766;
  wire [0:0] s_2767;
  wire [0:0] s_2768;
  wire [0:0] s_2769;
  wire [1:0] s_2770;
  wire [0:0] s_2771;
  wire [0:0] s_2772;
  wire [0:0] s_2773;
  wire [0:0] s_2774;
  wire [0:0] s_2775;
  wire [2:0] s_2776;
  wire [0:0] s_2777;
  wire [0:0] s_2778;
  wire [1:0] s_2779;
  wire [1:0] s_2780;
  wire [1:0] s_2781;
  wire [3:0] s_2782;
  wire [0:0] s_2783;
  wire [0:0] s_2784;
  wire [2:0] s_2785;
  wire [2:0] s_2786;
  wire [2:0] s_2787;
  wire [4:0] s_2788;
  wire [0:0] s_2789;
  wire [0:0] s_2790;
  wire [3:0] s_2791;
  wire [3:0] s_2792;
  wire [3:0] s_2793;
  wire [0:0] s_2794;
  wire [5:0] s_2795;
  wire [0:0] s_2796;
  wire [0:0] s_2797;
  wire [4:0] s_2798;
  wire [0:0] s_2799;
  wire [0:0] s_2800;
  wire [3:0] s_2801;
  wire [0:0] s_2802;
  wire [0:0] s_2803;
  wire [2:0] s_2804;
  wire [0:0] s_2805;
  wire [0:0] s_2806;
  wire [1:0] s_2807;
  wire [0:0] s_2808;
  wire [0:0] s_2809;
  wire [0:0] s_2810;
  wire [1:0] s_2811;
  wire [3:0] s_2812;
  wire [7:0] s_2813;
  wire [15:0] s_2814;
  wire [31:0] s_2815;
  wire [0:0] s_2816;
  wire [0:0] s_2817;
  wire [0:0] s_2818;
  wire [0:0] s_2819;
  wire [0:0] s_2820;
  wire [0:0] s_2821;
  wire [0:0] s_2822;
  wire [1:0] s_2823;
  wire [0:0] s_2824;
  wire [0:0] s_2825;
  wire [0:0] s_2826;
  wire [1:0] s_2827;
  wire [0:0] s_2828;
  wire [0:0] s_2829;
  wire [0:0] s_2830;
  wire [0:0] s_2831;
  wire [0:0] s_2832;
  wire [0:0] s_2833;
  wire [1:0] s_2834;
  wire [0:0] s_2835;
  wire [0:0] s_2836;
  wire [0:0] s_2837;
  wire [0:0] s_2838;
  wire [0:0] s_2839;
  wire [0:0] s_2840;
  wire [2:0] s_2841;
  wire [0:0] s_2842;
  wire [0:0] s_2843;
  wire [1:0] s_2844;
  wire [0:0] s_2845;
  wire [0:0] s_2846;
  wire [0:0] s_2847;
  wire [1:0] s_2848;
  wire [3:0] s_2849;
  wire [0:0] s_2850;
  wire [0:0] s_2851;
  wire [0:0] s_2852;
  wire [0:0] s_2853;
  wire [0:0] s_2854;
  wire [0:0] s_2855;
  wire [0:0] s_2856;
  wire [1:0] s_2857;
  wire [0:0] s_2858;
  wire [0:0] s_2859;
  wire [0:0] s_2860;
  wire [1:0] s_2861;
  wire [0:0] s_2862;
  wire [0:0] s_2863;
  wire [0:0] s_2864;
  wire [0:0] s_2865;
  wire [0:0] s_2866;
  wire [0:0] s_2867;
  wire [1:0] s_2868;
  wire [0:0] s_2869;
  wire [0:0] s_2870;
  wire [0:0] s_2871;
  wire [0:0] s_2872;
  wire [0:0] s_2873;
  wire [2:0] s_2874;
  wire [0:0] s_2875;
  wire [0:0] s_2876;
  wire [1:0] s_2877;
  wire [1:0] s_2878;
  wire [1:0] s_2879;
  wire [0:0] s_2880;
  wire [3:0] s_2881;
  wire [0:0] s_2882;
  wire [0:0] s_2883;
  wire [2:0] s_2884;
  wire [0:0] s_2885;
  wire [0:0] s_2886;
  wire [1:0] s_2887;
  wire [0:0] s_2888;
  wire [0:0] s_2889;
  wire [0:0] s_2890;
  wire [1:0] s_2891;
  wire [3:0] s_2892;
  wire [7:0] s_2893;
  wire [0:0] s_2894;
  wire [0:0] s_2895;
  wire [0:0] s_2896;
  wire [0:0] s_2897;
  wire [0:0] s_2898;
  wire [0:0] s_2899;
  wire [0:0] s_2900;
  wire [1:0] s_2901;
  wire [0:0] s_2902;
  wire [0:0] s_2903;
  wire [0:0] s_2904;
  wire [1:0] s_2905;
  wire [0:0] s_2906;
  wire [0:0] s_2907;
  wire [0:0] s_2908;
  wire [0:0] s_2909;
  wire [0:0] s_2910;
  wire [0:0] s_2911;
  wire [1:0] s_2912;
  wire [0:0] s_2913;
  wire [0:0] s_2914;
  wire [0:0] s_2915;
  wire [0:0] s_2916;
  wire [0:0] s_2917;
  wire [0:0] s_2918;
  wire [2:0] s_2919;
  wire [0:0] s_2920;
  wire [0:0] s_2921;
  wire [1:0] s_2922;
  wire [0:0] s_2923;
  wire [0:0] s_2924;
  wire [0:0] s_2925;
  wire [1:0] s_2926;
  wire [3:0] s_2927;
  wire [0:0] s_2928;
  wire [0:0] s_2929;
  wire [0:0] s_2930;
  wire [0:0] s_2931;
  wire [0:0] s_2932;
  wire [0:0] s_2933;
  wire [0:0] s_2934;
  wire [1:0] s_2935;
  wire [0:0] s_2936;
  wire [0:0] s_2937;
  wire [0:0] s_2938;
  wire [1:0] s_2939;
  wire [0:0] s_2940;
  wire [0:0] s_2941;
  wire [0:0] s_2942;
  wire [0:0] s_2943;
  wire [0:0] s_2944;
  wire [0:0] s_2945;
  wire [1:0] s_2946;
  wire [0:0] s_2947;
  wire [0:0] s_2948;
  wire [0:0] s_2949;
  wire [0:0] s_2950;
  wire [0:0] s_2951;
  wire [2:0] s_2952;
  wire [0:0] s_2953;
  wire [0:0] s_2954;
  wire [1:0] s_2955;
  wire [1:0] s_2956;
  wire [1:0] s_2957;
  wire [3:0] s_2958;
  wire [0:0] s_2959;
  wire [0:0] s_2960;
  wire [2:0] s_2961;
  wire [2:0] s_2962;
  wire [2:0] s_2963;
  wire [0:0] s_2964;
  wire [4:0] s_2965;
  wire [0:0] s_2966;
  wire [0:0] s_2967;
  wire [3:0] s_2968;
  wire [0:0] s_2969;
  wire [0:0] s_2970;
  wire [2:0] s_2971;
  wire [0:0] s_2972;
  wire [0:0] s_2973;
  wire [1:0] s_2974;
  wire [0:0] s_2975;
  wire [0:0] s_2976;
  wire [0:0] s_2977;
  wire [1:0] s_2978;
  wire [3:0] s_2979;
  wire [7:0] s_2980;
  wire [15:0] s_2981;
  wire [0:0] s_2982;
  wire [0:0] s_2983;
  wire [0:0] s_2984;
  wire [0:0] s_2985;
  wire [0:0] s_2986;
  wire [0:0] s_2987;
  wire [0:0] s_2988;
  wire [1:0] s_2989;
  wire [0:0] s_2990;
  wire [0:0] s_2991;
  wire [0:0] s_2992;
  wire [1:0] s_2993;
  wire [0:0] s_2994;
  wire [0:0] s_2995;
  wire [0:0] s_2996;
  wire [0:0] s_2997;
  wire [0:0] s_2998;
  wire [0:0] s_2999;
  wire [1:0] s_3000;
  wire [0:0] s_3001;
  wire [0:0] s_3002;
  wire [0:0] s_3003;
  wire [0:0] s_3004;
  wire [0:0] s_3005;
  wire [0:0] s_3006;
  wire [2:0] s_3007;
  wire [0:0] s_3008;
  wire [0:0] s_3009;
  wire [1:0] s_3010;
  wire [0:0] s_3011;
  wire [0:0] s_3012;
  wire [0:0] s_3013;
  wire [1:0] s_3014;
  wire [3:0] s_3015;
  wire [0:0] s_3016;
  wire [0:0] s_3017;
  wire [0:0] s_3018;
  wire [0:0] s_3019;
  wire [0:0] s_3020;
  wire [0:0] s_3021;
  wire [0:0] s_3022;
  wire [1:0] s_3023;
  wire [0:0] s_3024;
  wire [0:0] s_3025;
  wire [0:0] s_3026;
  wire [1:0] s_3027;
  wire [0:0] s_3028;
  wire [0:0] s_3029;
  wire [0:0] s_3030;
  wire [0:0] s_3031;
  wire [0:0] s_3032;
  wire [0:0] s_3033;
  wire [1:0] s_3034;
  wire [0:0] s_3035;
  wire [0:0] s_3036;
  wire [0:0] s_3037;
  wire [0:0] s_3038;
  wire [0:0] s_3039;
  wire [2:0] s_3040;
  wire [0:0] s_3041;
  wire [0:0] s_3042;
  wire [1:0] s_3043;
  wire [1:0] s_3044;
  wire [1:0] s_3045;
  wire [0:0] s_3046;
  wire [3:0] s_3047;
  wire [0:0] s_3048;
  wire [0:0] s_3049;
  wire [2:0] s_3050;
  wire [0:0] s_3051;
  wire [0:0] s_3052;
  wire [1:0] s_3053;
  wire [0:0] s_3054;
  wire [0:0] s_3055;
  wire [0:0] s_3056;
  wire [1:0] s_3057;
  wire [3:0] s_3058;
  wire [7:0] s_3059;
  wire [0:0] s_3060;
  wire [0:0] s_3061;
  wire [0:0] s_3062;
  wire [0:0] s_3063;
  wire [0:0] s_3064;
  wire [0:0] s_3065;
  wire [0:0] s_3066;
  wire [1:0] s_3067;
  wire [0:0] s_3068;
  wire [0:0] s_3069;
  wire [0:0] s_3070;
  wire [1:0] s_3071;
  wire [0:0] s_3072;
  wire [0:0] s_3073;
  wire [0:0] s_3074;
  wire [0:0] s_3075;
  wire [0:0] s_3076;
  wire [0:0] s_3077;
  wire [1:0] s_3078;
  wire [0:0] s_3079;
  wire [0:0] s_3080;
  wire [0:0] s_3081;
  wire [0:0] s_3082;
  wire [0:0] s_3083;
  wire [0:0] s_3084;
  wire [2:0] s_3085;
  wire [0:0] s_3086;
  wire [0:0] s_3087;
  wire [1:0] s_3088;
  wire [0:0] s_3089;
  wire [0:0] s_3090;
  wire [0:0] s_3091;
  wire [1:0] s_3092;
  wire [3:0] s_3093;
  wire [0:0] s_3094;
  wire [0:0] s_3095;
  wire [0:0] s_3096;
  wire [0:0] s_3097;
  wire [0:0] s_3098;
  wire [0:0] s_3099;
  wire [0:0] s_3100;
  wire [1:0] s_3101;
  wire [0:0] s_3102;
  wire [0:0] s_3103;
  wire [0:0] s_3104;
  wire [1:0] s_3105;
  wire [0:0] s_3106;
  wire [0:0] s_3107;
  wire [0:0] s_3108;
  wire [0:0] s_3109;
  wire [0:0] s_3110;
  wire [0:0] s_3111;
  wire [1:0] s_3112;
  wire [0:0] s_3113;
  wire [0:0] s_3114;
  wire [0:0] s_3115;
  wire [0:0] s_3116;
  wire [0:0] s_3117;
  wire [2:0] s_3118;
  wire [0:0] s_3119;
  wire [0:0] s_3120;
  wire [1:0] s_3121;
  wire [1:0] s_3122;
  wire [1:0] s_3123;
  wire [3:0] s_3124;
  wire [0:0] s_3125;
  wire [0:0] s_3126;
  wire [2:0] s_3127;
  wire [2:0] s_3128;
  wire [2:0] s_3129;
  wire [4:0] s_3130;
  wire [0:0] s_3131;
  wire [0:0] s_3132;
  wire [3:0] s_3133;
  wire [3:0] s_3134;
  wire [3:0] s_3135;
  wire [5:0] s_3136;
  wire [0:0] s_3137;
  wire [0:0] s_3138;
  wire [4:0] s_3139;
  wire [4:0] s_3140;
  wire [4:0] s_3141;
  wire [12:0] s_3142;
  wire [12:0] s_3143;
  wire [12:0] s_3144;
  wire [12:0] s_3145;
  wire [12:0] s_3146;
  wire [12:0] s_3147;
  wire [0:0] s_3148;
  wire [12:0] s_3149;
  wire [12:0] s_3150;
  wire [1:0] s_3151;
  wire [0:0] s_3152;
  wire [52:0] s_3153;
  wire [0:0] s_3154;
  wire [0:0] s_3155;
  wire [0:0] s_3156;
  wire [0:0] s_3157;
  wire [0:0] s_3158;
  wire [0:0] s_3159;
  wire [0:0] s_3160;
  wire [0:0] s_3161;
  wire [0:0] s_3162;
  wire [0:0] s_3163;
  wire [0:0] s_3164;
  wire [0:0] s_3165;
  wire [56:0] s_3166;
  wire [56:0] s_3167;
  wire [0:0] s_3168;
  wire [0:0] s_3169;
  wire [0:0] s_3170;
  wire [52:0] s_3171;
  wire [0:0] s_3172;
  wire [0:0] s_3173;
  wire [0:0] s_3174;
  wire [0:0] s_3175;
  wire [10:0] s_3176;
  wire [0:0] s_3177;
  wire [51:0] s_3178;
  wire [63:0] s_3179;
  wire [11:0] s_3180;
  wire [0:0] s_3181;
  wire [10:0] s_3182;
  wire [10:0] s_3183;
  wire [12:0] s_3184;
  wire [12:0] s_3185;
  wire [12:0] s_3186;
  wire [12:0] s_3187;
  wire [12:0] s_3188;
  wire [12:0] s_3189;
  wire [9:0] s_3190;
  wire [51:0] s_3191;
  wire [0:0] s_3192;
  wire [0:0] s_3193;
  wire [10:0] s_3194;
  wire [0:0] s_3195;
  wire [0:0] s_3196;
  wire [0:0] s_3197;
  wire [52:0] s_3198;
  wire [0:0] s_3199;
  wire [0:0] s_3200;
  wire [0:0] s_3201;
  wire [0:0] s_3202;
  wire [0:0] s_3203;
  wire [11:0] s_3204;
  wire [0:0] s_3205;
  wire [0:0] s_3206;
  wire [0:0] s_3207;
  wire [10:0] s_3208;
  wire [0:0] s_3209;
  wire [51:0] s_3210;
  wire [0:0] s_3211;
  wire [0:0] s_3212;
  wire [0:0] s_3213;
  wire [0:0] s_3214;
  wire [0:0] s_3215;
  wire [0:0] s_3216;
  wire [0:0] s_3217;
  wire [0:0] s_3218;
  wire [0:0] s_3219;
  wire [0:0] s_3220;
  wire [10:0] s_3221;
  wire [0:0] s_3222;
  wire [51:0] s_3223;
  wire [0:0] s_3224;
  wire [0:0] s_3225;
  wire [10:0] s_3226;
  wire [0:0] s_3227;
  wire [51:0] s_3228;
  wire [0:0] s_3229;

  assign s_0 = s_3216?s_1:s_9;
  dq #(64, 65) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_8};
  assign s_3 = s_4 ^ s_6;
  assign s_4 = s_5[63];
  assign s_5 = double_div_a;
  assign s_6 = s_7[63];
  assign s_7 = double_div_b;
  assign s_8 = 63'd9221120237041090560;
  assign s_9 = s_3199?s_10:s_13;
  dq #(64, 65) dq_s_10 (clk, s_10, s_11);
  assign s_11 = {s_3,s_12};
  assign s_12 = 63'd9218868437227405312;
  assign s_13 = s_3197?s_14:s_17;
  dq #(64, 65) dq_s_14 (clk, s_14, s_15);
  assign s_15 = {s_3,s_16};
  assign s_16 = 63'd0;
  assign s_17 = s_3192?s_18:s_3179;
  assign s_18 = {s_19,s_22};
  dq #(12, 65) dq_s_19 (clk, s_19, s_20);
  assign s_20 = {s_3,s_21};
  assign s_21 = 11'd0;
  assign s_22 = s_23[51:0];
  assign s_23 = s_3173?s_24:s_25;
  assign s_24 = 1'd0;
  dq #(53, 1) dq_s_25 (clk, s_25, s_26);
  assign s_26 = s_3172?s_27:s_3171;
  assign s_27 = s_28[53:1];
  assign s_28 = s_3154?s_29:s_3153;
  dq #(54, 1) dq_s_29 (clk, s_29, s_30);
  assign s_30 = s_31 + s_3152;
  assign s_31 = s_32;
  assign s_32 = s_33[52:0];
  assign s_33 = s_34 >> s_3151;
  dq #(56, 1) dq_s_34 (clk, s_34, s_35);
  assign s_35 = s_36 << s_2431;
  dq #(56, 2) dq_s_36 (clk, s_36, s_37);
  dq #(56, 1) dq_s_37 (clk, s_37, s_38);
  assign s_38 = s_39 >> s_2415;
  dq #(56, 1) dq_s_39 (clk, s_39, s_40);
  assign s_40 = s_2405?s_41:s_2403;
  assign s_41 = s_42 << s_2402;
  dq #(56, 1) dq_s_42 (clk, s_42, s_43);
  assign s_43 = s_2392?s_44:s_2390;
  assign s_44 = s_45 << s_2389;
  dq #(56, 1) dq_s_45 (clk, s_45, s_46);
  assign s_46 = s_2379?s_47:s_2377;
  assign s_47 = s_48 << s_2376;
  dq #(56, 1) dq_s_48 (clk, s_48, s_49);
  assign s_49 = s_2366?s_50:s_2364;
  assign s_50 = s_51 << s_2363;
  dq #(56, 1) dq_s_51 (clk, s_51, s_52);
  assign s_52 = s_2353?s_53:s_2351;
  assign s_53 = s_54 << s_2350;
  dq #(56, 1) dq_s_54 (clk, s_54, s_55);
  assign s_55 = s_2340?s_56:s_2338;
  assign s_56 = s_57 << s_2337;
  dq #(56, 1) dq_s_57 (clk, s_57, s_58);
  assign s_58 = s_2327?s_59:s_2325;
  assign s_59 = s_60 << s_2324;
  dq #(56, 1) dq_s_60 (clk, s_60, s_61);
  assign s_61 = s_2314?s_62:s_2312;
  assign s_62 = s_63 << s_2311;
  dq #(56, 1) dq_s_63 (clk, s_63, s_64);
  assign s_64 = s_2301?s_65:s_2299;
  assign s_65 = s_66 << s_2298;
  dq #(56, 1) dq_s_66 (clk, s_66, s_67);
  assign s_67 = s_2288?s_68:s_2286;
  assign s_68 = s_69 << s_2285;
  dq #(56, 1) dq_s_69 (clk, s_69, s_70);
  assign s_70 = s_2275?s_71:s_2273;
  assign s_71 = s_72 << s_2272;
  dq #(56, 1) dq_s_72 (clk, s_72, s_73);
  assign s_73 = s_2262?s_74:s_2260;
  assign s_74 = s_75 << s_2259;
  dq #(56, 1) dq_s_75 (clk, s_75, s_76);
  assign s_76 = s_2249?s_77:s_2247;
  assign s_77 = s_78 << s_2246;
  dq #(56, 1) dq_s_78 (clk, s_78, s_79);
  assign s_79 = s_2236?s_80:s_2234;
  assign s_80 = s_81 << s_2233;
  dq #(56, 1) dq_s_81 (clk, s_81, s_82);
  assign s_82 = s_2223?s_83:s_2221;
  assign s_83 = s_84 << s_2220;
  dq #(56, 1) dq_s_84 (clk, s_84, s_85);
  assign s_85 = s_2210?s_86:s_2208;
  assign s_86 = s_87 << s_2207;
  dq #(56, 1) dq_s_87 (clk, s_87, s_88);
  assign s_88 = s_2197?s_89:s_2195;
  assign s_89 = s_90 << s_2194;
  dq #(56, 1) dq_s_90 (clk, s_90, s_91);
  assign s_91 = s_2184?s_92:s_2182;
  assign s_92 = s_93 << s_2181;
  dq #(56, 1) dq_s_93 (clk, s_93, s_94);
  assign s_94 = s_2171?s_95:s_2169;
  assign s_95 = s_96 << s_2168;
  dq #(56, 1) dq_s_96 (clk, s_96, s_97);
  assign s_97 = s_2158?s_98:s_2156;
  assign s_98 = s_99 << s_2155;
  dq #(56, 1) dq_s_99 (clk, s_99, s_100);
  assign s_100 = s_2145?s_101:s_2143;
  assign s_101 = s_102 << s_2142;
  dq #(56, 1) dq_s_102 (clk, s_102, s_103);
  assign s_103 = s_2132?s_104:s_2130;
  assign s_104 = s_105 << s_2129;
  dq #(56, 1) dq_s_105 (clk, s_105, s_106);
  assign s_106 = s_2119?s_107:s_2117;
  assign s_107 = s_108 << s_2116;
  dq #(56, 1) dq_s_108 (clk, s_108, s_109);
  assign s_109 = s_2106?s_110:s_2104;
  assign s_110 = s_111 << s_2103;
  dq #(56, 1) dq_s_111 (clk, s_111, s_112);
  assign s_112 = s_2093?s_113:s_2091;
  assign s_113 = s_114 << s_2090;
  dq #(56, 1) dq_s_114 (clk, s_114, s_115);
  assign s_115 = s_2080?s_116:s_2078;
  assign s_116 = s_117 << s_2077;
  dq #(56, 1) dq_s_117 (clk, s_117, s_118);
  assign s_118 = s_2067?s_119:s_2065;
  assign s_119 = s_120 << s_2064;
  dq #(56, 1) dq_s_120 (clk, s_120, s_121);
  assign s_121 = s_2054?s_122:s_2052;
  assign s_122 = s_123 << s_2051;
  dq #(56, 1) dq_s_123 (clk, s_123, s_124);
  assign s_124 = s_2041?s_125:s_2039;
  assign s_125 = s_126 << s_2038;
  dq #(56, 1) dq_s_126 (clk, s_126, s_127);
  assign s_127 = s_2028?s_128:s_2026;
  assign s_128 = s_129 << s_2025;
  dq #(56, 1) dq_s_129 (clk, s_129, s_130);
  assign s_130 = s_2015?s_131:s_2013;
  assign s_131 = s_132 << s_2012;
  dq #(56, 1) dq_s_132 (clk, s_132, s_133);
  assign s_133 = s_2002?s_134:s_2000;
  assign s_134 = s_135 << s_1999;
  dq #(56, 1) dq_s_135 (clk, s_135, s_136);
  assign s_136 = s_1989?s_137:s_1987;
  assign s_137 = s_138 << s_1986;
  dq #(56, 1) dq_s_138 (clk, s_138, s_139);
  assign s_139 = s_1976?s_140:s_1974;
  assign s_140 = s_141 << s_1973;
  dq #(56, 1) dq_s_141 (clk, s_141, s_142);
  assign s_142 = s_1963?s_143:s_1961;
  assign s_143 = s_144 << s_1960;
  dq #(56, 1) dq_s_144 (clk, s_144, s_145);
  assign s_145 = s_1950?s_146:s_1948;
  assign s_146 = s_147 << s_1947;
  dq #(56, 1) dq_s_147 (clk, s_147, s_148);
  assign s_148 = s_1937?s_149:s_1935;
  assign s_149 = s_150 << s_1934;
  dq #(56, 1) dq_s_150 (clk, s_150, s_151);
  assign s_151 = s_1924?s_152:s_1922;
  assign s_152 = s_153 << s_1921;
  dq #(56, 1) dq_s_153 (clk, s_153, s_154);
  assign s_154 = s_1911?s_155:s_1909;
  assign s_155 = s_156 << s_1908;
  dq #(56, 1) dq_s_156 (clk, s_156, s_157);
  assign s_157 = s_1898?s_158:s_1896;
  assign s_158 = s_159 << s_1895;
  dq #(56, 1) dq_s_159 (clk, s_159, s_160);
  assign s_160 = s_1885?s_161:s_1883;
  assign s_161 = s_162 << s_1882;
  dq #(56, 1) dq_s_162 (clk, s_162, s_163);
  assign s_163 = s_1872?s_164:s_1870;
  assign s_164 = s_165 << s_1869;
  dq #(56, 1) dq_s_165 (clk, s_165, s_166);
  assign s_166 = s_1859?s_167:s_1857;
  assign s_167 = s_168 << s_1856;
  dq #(56, 1) dq_s_168 (clk, s_168, s_169);
  assign s_169 = s_1846?s_170:s_1844;
  assign s_170 = s_171 << s_1843;
  dq #(56, 1) dq_s_171 (clk, s_171, s_172);
  assign s_172 = s_1833?s_173:s_1831;
  assign s_173 = s_174 << s_1830;
  dq #(56, 1) dq_s_174 (clk, s_174, s_175);
  assign s_175 = s_1820?s_176:s_1818;
  assign s_176 = s_177 << s_1817;
  dq #(56, 1) dq_s_177 (clk, s_177, s_178);
  assign s_178 = s_1807?s_179:s_1805;
  assign s_179 = s_180 << s_1804;
  dq #(56, 1) dq_s_180 (clk, s_180, s_181);
  assign s_181 = s_1794?s_182:s_1792;
  assign s_182 = s_183 << s_1791;
  dq #(56, 1) dq_s_183 (clk, s_183, s_184);
  assign s_184 = s_1781?s_185:s_1779;
  assign s_185 = s_186 << s_1778;
  dq #(56, 1) dq_s_186 (clk, s_186, s_187);
  assign s_187 = s_1768?s_188:s_1766;
  assign s_188 = s_189 << s_1765;
  dq #(56, 1) dq_s_189 (clk, s_189, s_190);
  assign s_190 = s_1755?s_191:s_1753;
  assign s_191 = s_192 << s_1752;
  dq #(56, 1) dq_s_192 (clk, s_192, s_193);
  assign s_193 = s_1742?s_194:s_1740;
  assign s_194 = s_195 << s_1739;
  dq #(56, 1) dq_s_195 (clk, s_195, s_196);
  assign s_196 = s_1729?s_197:s_1727;
  assign s_197 = s_198 << s_1726;
  dq #(56, 1) dq_s_198 (clk, s_198, s_199);
  assign s_199 = s_1716?s_200:s_1714;
  assign s_200 = s_201 << s_1713;
  dq #(56, 1) dq_s_201 (clk, s_201, s_202);
  assign s_202 = s_1703?s_203:s_1701;
  assign s_203 = s_204 << s_1700;
  dq #(56, 1) dq_s_204 (clk, s_204, s_205);
  assign s_205 = s_213?s_206:s_210;
  dq #(56, 3) dq_s_206 (clk, s_206, s_207);
  assign s_207 = s_208 << s_209;
  assign s_208 = 56'd0;
  assign s_209 = 1'd1;
  dq #(56, 3) dq_s_210 (clk, s_210, s_211);
  assign s_211 = s_207 | s_212;
  assign s_212 = 1'd1;
  assign s_213 = s_214[56];
  assign s_214 = s_215 - s_958;
  assign s_215 = s_216;
  assign s_216 = s_217 << s_957;
  assign s_217 = s_218;
  dq #(53, 1) dq_s_218 (clk, s_218, s_219);
  assign s_219 = s_220 << s_231;
  dq #(53, 2) dq_s_220 (clk, s_220, s_221);
  assign s_221 = {s_222,s_230};
  assign s_222 = s_225?s_223:s_224;
  assign s_223 = 1'd0;
  assign s_224 = 1'd1;
  assign s_225 = s_226 == s_229;
  assign s_226 = s_227 - s_228;
  assign s_227 = s_5[62:52];
  assign s_228 = 10'd1023;
  assign s_229 = -11'd1023;
  assign s_230 = s_5[51:0];
  dq #(13, 1) dq_s_231 (clk, s_231, s_232);
  assign s_232 = s_954?s_233:s_948;
  dq #(7, 1) dq_s_233 (clk, s_233, s_234);
  assign s_234 = {s_235,s_942};
  assign s_235 = s_236 & s_600;
  assign s_236 = s_237[5];
  assign s_237 = {s_238,s_594};
  assign s_238 = s_239 & s_428;
  assign s_239 = s_240[4];
  assign s_240 = {s_241,s_422};
  assign s_241 = s_242 & s_344;
  assign s_242 = s_243[3];
  assign s_243 = {s_244,s_338};
  assign s_244 = s_245 & s_304;
  assign s_245 = s_246[2];
  assign s_246 = {s_247,s_298};
  assign s_247 = s_248 & s_286;
  assign s_248 = s_249[1];
  assign s_249 = {s_250,s_282};
  assign s_250 = s_251 & s_280;
  assign s_251 = ~s_252;
  assign s_252 = s_253[1];
  assign s_253 = s_254[3:2];
  assign s_254 = s_255[7:4];
  assign s_255 = s_256[15:8];
  assign s_256 = s_257[31:16];
  assign s_257 = s_258[63:32];
  assign s_258 = {s_259,s_279};
  assign s_259 = {s_260,s_278};
  assign s_260 = {s_261,s_277};
  assign s_261 = {s_262,s_276};
  assign s_262 = {s_263,s_275};
  assign s_263 = {s_264,s_274};
  assign s_264 = {s_265,s_273};
  assign s_265 = {s_266,s_272};
  assign s_266 = {s_267,s_271};
  assign s_267 = {s_268,s_270};
  assign s_268 = {s_221,s_269};
  assign s_269 = 1'd1;
  assign s_270 = 1'd1;
  assign s_271 = 1'd1;
  assign s_272 = 1'd1;
  assign s_273 = 1'd1;
  assign s_274 = 1'd1;
  assign s_275 = 1'd1;
  assign s_276 = 1'd1;
  assign s_277 = 1'd1;
  assign s_278 = 1'd1;
  assign s_279 = 1'd1;
  assign s_280 = ~s_281;
  assign s_281 = s_253[0];
  assign s_282 = s_283 & s_285;
  assign s_283 = ~s_284;
  assign s_284 = s_253[1];
  assign s_285 = s_253[0];
  assign s_286 = s_287[1];
  assign s_287 = {s_288,s_294};
  assign s_288 = s_289 & s_292;
  assign s_289 = ~s_290;
  assign s_290 = s_291[1];
  assign s_291 = s_254[1:0];
  assign s_292 = ~s_293;
  assign s_293 = s_291[0];
  assign s_294 = s_295 & s_297;
  assign s_295 = ~s_296;
  assign s_296 = s_291[1];
  assign s_297 = s_291[0];
  assign s_298 = {s_299,s_301};
  assign s_299 = s_248 & s_300;
  assign s_300 = ~s_286;
  assign s_301 = s_248?s_302:s_303;
  assign s_302 = s_287[0:0];
  assign s_303 = s_249[0:0];
  assign s_304 = s_305[2];
  assign s_305 = {s_306,s_332};
  assign s_306 = s_307 & s_320;
  assign s_307 = s_308[1];
  assign s_308 = {s_309,s_316};
  assign s_309 = s_310 & s_314;
  assign s_310 = ~s_311;
  assign s_311 = s_312[1];
  assign s_312 = s_313[3:2];
  assign s_313 = s_255[3:0];
  assign s_314 = ~s_315;
  assign s_315 = s_312[0];
  assign s_316 = s_317 & s_319;
  assign s_317 = ~s_318;
  assign s_318 = s_312[1];
  assign s_319 = s_312[0];
  assign s_320 = s_321[1];
  assign s_321 = {s_322,s_328};
  assign s_322 = s_323 & s_326;
  assign s_323 = ~s_324;
  assign s_324 = s_325[1];
  assign s_325 = s_313[1:0];
  assign s_326 = ~s_327;
  assign s_327 = s_325[0];
  assign s_328 = s_329 & s_331;
  assign s_329 = ~s_330;
  assign s_330 = s_325[1];
  assign s_331 = s_325[0];
  assign s_332 = {s_333,s_335};
  assign s_333 = s_307 & s_334;
  assign s_334 = ~s_320;
  assign s_335 = s_307?s_336:s_337;
  assign s_336 = s_321[0:0];
  assign s_337 = s_308[0:0];
  assign s_338 = {s_339,s_341};
  assign s_339 = s_245 & s_340;
  assign s_340 = ~s_304;
  assign s_341 = s_245?s_342:s_343;
  assign s_342 = s_305[1:0];
  assign s_343 = s_246[1:0];
  assign s_344 = s_345[3];
  assign s_345 = {s_346,s_416};
  assign s_346 = s_347 & s_382;
  assign s_347 = s_348[2];
  assign s_348 = {s_349,s_376};
  assign s_349 = s_350 & s_364;
  assign s_350 = s_351[1];
  assign s_351 = {s_352,s_360};
  assign s_352 = s_353 & s_358;
  assign s_353 = ~s_354;
  assign s_354 = s_355[1];
  assign s_355 = s_356[3:2];
  assign s_356 = s_357[7:4];
  assign s_357 = s_256[7:0];
  assign s_358 = ~s_359;
  assign s_359 = s_355[0];
  assign s_360 = s_361 & s_363;
  assign s_361 = ~s_362;
  assign s_362 = s_355[1];
  assign s_363 = s_355[0];
  assign s_364 = s_365[1];
  assign s_365 = {s_366,s_372};
  assign s_366 = s_367 & s_370;
  assign s_367 = ~s_368;
  assign s_368 = s_369[1];
  assign s_369 = s_356[1:0];
  assign s_370 = ~s_371;
  assign s_371 = s_369[0];
  assign s_372 = s_373 & s_375;
  assign s_373 = ~s_374;
  assign s_374 = s_369[1];
  assign s_375 = s_369[0];
  assign s_376 = {s_377,s_379};
  assign s_377 = s_350 & s_378;
  assign s_378 = ~s_364;
  assign s_379 = s_350?s_380:s_381;
  assign s_380 = s_365[0:0];
  assign s_381 = s_351[0:0];
  assign s_382 = s_383[2];
  assign s_383 = {s_384,s_410};
  assign s_384 = s_385 & s_398;
  assign s_385 = s_386[1];
  assign s_386 = {s_387,s_394};
  assign s_387 = s_388 & s_392;
  assign s_388 = ~s_389;
  assign s_389 = s_390[1];
  assign s_390 = s_391[3:2];
  assign s_391 = s_357[3:0];
  assign s_392 = ~s_393;
  assign s_393 = s_390[0];
  assign s_394 = s_395 & s_397;
  assign s_395 = ~s_396;
  assign s_396 = s_390[1];
  assign s_397 = s_390[0];
  assign s_398 = s_399[1];
  assign s_399 = {s_400,s_406};
  assign s_400 = s_401 & s_404;
  assign s_401 = ~s_402;
  assign s_402 = s_403[1];
  assign s_403 = s_391[1:0];
  assign s_404 = ~s_405;
  assign s_405 = s_403[0];
  assign s_406 = s_407 & s_409;
  assign s_407 = ~s_408;
  assign s_408 = s_403[1];
  assign s_409 = s_403[0];
  assign s_410 = {s_411,s_413};
  assign s_411 = s_385 & s_412;
  assign s_412 = ~s_398;
  assign s_413 = s_385?s_414:s_415;
  assign s_414 = s_399[0:0];
  assign s_415 = s_386[0:0];
  assign s_416 = {s_417,s_419};
  assign s_417 = s_347 & s_418;
  assign s_418 = ~s_382;
  assign s_419 = s_347?s_420:s_421;
  assign s_420 = s_383[1:0];
  assign s_421 = s_348[1:0];
  assign s_422 = {s_423,s_425};
  assign s_423 = s_242 & s_424;
  assign s_424 = ~s_344;
  assign s_425 = s_242?s_426:s_427;
  assign s_426 = s_345[2:0];
  assign s_427 = s_243[2:0];
  assign s_428 = s_429[4];
  assign s_429 = {s_430,s_588};
  assign s_430 = s_431 & s_510;
  assign s_431 = s_432[3];
  assign s_432 = {s_433,s_504};
  assign s_433 = s_434 & s_470;
  assign s_434 = s_435[2];
  assign s_435 = {s_436,s_464};
  assign s_436 = s_437 & s_452;
  assign s_437 = s_438[1];
  assign s_438 = {s_439,s_448};
  assign s_439 = s_440 & s_446;
  assign s_440 = ~s_441;
  assign s_441 = s_442[1];
  assign s_442 = s_443[3:2];
  assign s_443 = s_444[7:4];
  assign s_444 = s_445[15:8];
  assign s_445 = s_257[15:0];
  assign s_446 = ~s_447;
  assign s_447 = s_442[0];
  assign s_448 = s_449 & s_451;
  assign s_449 = ~s_450;
  assign s_450 = s_442[1];
  assign s_451 = s_442[0];
  assign s_452 = s_453[1];
  assign s_453 = {s_454,s_460};
  assign s_454 = s_455 & s_458;
  assign s_455 = ~s_456;
  assign s_456 = s_457[1];
  assign s_457 = s_443[1:0];
  assign s_458 = ~s_459;
  assign s_459 = s_457[0];
  assign s_460 = s_461 & s_463;
  assign s_461 = ~s_462;
  assign s_462 = s_457[1];
  assign s_463 = s_457[0];
  assign s_464 = {s_465,s_467};
  assign s_465 = s_437 & s_466;
  assign s_466 = ~s_452;
  assign s_467 = s_437?s_468:s_469;
  assign s_468 = s_453[0:0];
  assign s_469 = s_438[0:0];
  assign s_470 = s_471[2];
  assign s_471 = {s_472,s_498};
  assign s_472 = s_473 & s_486;
  assign s_473 = s_474[1];
  assign s_474 = {s_475,s_482};
  assign s_475 = s_476 & s_480;
  assign s_476 = ~s_477;
  assign s_477 = s_478[1];
  assign s_478 = s_479[3:2];
  assign s_479 = s_444[3:0];
  assign s_480 = ~s_481;
  assign s_481 = s_478[0];
  assign s_482 = s_483 & s_485;
  assign s_483 = ~s_484;
  assign s_484 = s_478[1];
  assign s_485 = s_478[0];
  assign s_486 = s_487[1];
  assign s_487 = {s_488,s_494};
  assign s_488 = s_489 & s_492;
  assign s_489 = ~s_490;
  assign s_490 = s_491[1];
  assign s_491 = s_479[1:0];
  assign s_492 = ~s_493;
  assign s_493 = s_491[0];
  assign s_494 = s_495 & s_497;
  assign s_495 = ~s_496;
  assign s_496 = s_491[1];
  assign s_497 = s_491[0];
  assign s_498 = {s_499,s_501};
  assign s_499 = s_473 & s_500;
  assign s_500 = ~s_486;
  assign s_501 = s_473?s_502:s_503;
  assign s_502 = s_487[0:0];
  assign s_503 = s_474[0:0];
  assign s_504 = {s_505,s_507};
  assign s_505 = s_434 & s_506;
  assign s_506 = ~s_470;
  assign s_507 = s_434?s_508:s_509;
  assign s_508 = s_471[1:0];
  assign s_509 = s_435[1:0];
  assign s_510 = s_511[3];
  assign s_511 = {s_512,s_582};
  assign s_512 = s_513 & s_548;
  assign s_513 = s_514[2];
  assign s_514 = {s_515,s_542};
  assign s_515 = s_516 & s_530;
  assign s_516 = s_517[1];
  assign s_517 = {s_518,s_526};
  assign s_518 = s_519 & s_524;
  assign s_519 = ~s_520;
  assign s_520 = s_521[1];
  assign s_521 = s_522[3:2];
  assign s_522 = s_523[7:4];
  assign s_523 = s_445[7:0];
  assign s_524 = ~s_525;
  assign s_525 = s_521[0];
  assign s_526 = s_527 & s_529;
  assign s_527 = ~s_528;
  assign s_528 = s_521[1];
  assign s_529 = s_521[0];
  assign s_530 = s_531[1];
  assign s_531 = {s_532,s_538};
  assign s_532 = s_533 & s_536;
  assign s_533 = ~s_534;
  assign s_534 = s_535[1];
  assign s_535 = s_522[1:0];
  assign s_536 = ~s_537;
  assign s_537 = s_535[0];
  assign s_538 = s_539 & s_541;
  assign s_539 = ~s_540;
  assign s_540 = s_535[1];
  assign s_541 = s_535[0];
  assign s_542 = {s_543,s_545};
  assign s_543 = s_516 & s_544;
  assign s_544 = ~s_530;
  assign s_545 = s_516?s_546:s_547;
  assign s_546 = s_531[0:0];
  assign s_547 = s_517[0:0];
  assign s_548 = s_549[2];
  assign s_549 = {s_550,s_576};
  assign s_550 = s_551 & s_564;
  assign s_551 = s_552[1];
  assign s_552 = {s_553,s_560};
  assign s_553 = s_554 & s_558;
  assign s_554 = ~s_555;
  assign s_555 = s_556[1];
  assign s_556 = s_557[3:2];
  assign s_557 = s_523[3:0];
  assign s_558 = ~s_559;
  assign s_559 = s_556[0];
  assign s_560 = s_561 & s_563;
  assign s_561 = ~s_562;
  assign s_562 = s_556[1];
  assign s_563 = s_556[0];
  assign s_564 = s_565[1];
  assign s_565 = {s_566,s_572};
  assign s_566 = s_567 & s_570;
  assign s_567 = ~s_568;
  assign s_568 = s_569[1];
  assign s_569 = s_557[1:0];
  assign s_570 = ~s_571;
  assign s_571 = s_569[0];
  assign s_572 = s_573 & s_575;
  assign s_573 = ~s_574;
  assign s_574 = s_569[1];
  assign s_575 = s_569[0];
  assign s_576 = {s_577,s_579};
  assign s_577 = s_551 & s_578;
  assign s_578 = ~s_564;
  assign s_579 = s_551?s_580:s_581;
  assign s_580 = s_565[0:0];
  assign s_581 = s_552[0:0];
  assign s_582 = {s_583,s_585};
  assign s_583 = s_513 & s_584;
  assign s_584 = ~s_548;
  assign s_585 = s_513?s_586:s_587;
  assign s_586 = s_549[1:0];
  assign s_587 = s_514[1:0];
  assign s_588 = {s_589,s_591};
  assign s_589 = s_431 & s_590;
  assign s_590 = ~s_510;
  assign s_591 = s_431?s_592:s_593;
  assign s_592 = s_511[2:0];
  assign s_593 = s_432[2:0];
  assign s_594 = {s_595,s_597};
  assign s_595 = s_239 & s_596;
  assign s_596 = ~s_428;
  assign s_597 = s_239?s_598:s_599;
  assign s_598 = s_429[3:0];
  assign s_599 = s_240[3:0];
  assign s_600 = s_601[5];
  assign s_601 = {s_602,s_936};
  assign s_602 = s_603 & s_770;
  assign s_603 = s_604[4];
  assign s_604 = {s_605,s_764};
  assign s_605 = s_606 & s_686;
  assign s_606 = s_607[3];
  assign s_607 = {s_608,s_680};
  assign s_608 = s_609 & s_646;
  assign s_609 = s_610[2];
  assign s_610 = {s_611,s_640};
  assign s_611 = s_612 & s_628;
  assign s_612 = s_613[1];
  assign s_613 = {s_614,s_624};
  assign s_614 = s_615 & s_622;
  assign s_615 = ~s_616;
  assign s_616 = s_617[1];
  assign s_617 = s_618[3:2];
  assign s_618 = s_619[7:4];
  assign s_619 = s_620[15:8];
  assign s_620 = s_621[31:16];
  assign s_621 = s_258[31:0];
  assign s_622 = ~s_623;
  assign s_623 = s_617[0];
  assign s_624 = s_625 & s_627;
  assign s_625 = ~s_626;
  assign s_626 = s_617[1];
  assign s_627 = s_617[0];
  assign s_628 = s_629[1];
  assign s_629 = {s_630,s_636};
  assign s_630 = s_631 & s_634;
  assign s_631 = ~s_632;
  assign s_632 = s_633[1];
  assign s_633 = s_618[1:0];
  assign s_634 = ~s_635;
  assign s_635 = s_633[0];
  assign s_636 = s_637 & s_639;
  assign s_637 = ~s_638;
  assign s_638 = s_633[1];
  assign s_639 = s_633[0];
  assign s_640 = {s_641,s_643};
  assign s_641 = s_612 & s_642;
  assign s_642 = ~s_628;
  assign s_643 = s_612?s_644:s_645;
  assign s_644 = s_629[0:0];
  assign s_645 = s_613[0:0];
  assign s_646 = s_647[2];
  assign s_647 = {s_648,s_674};
  assign s_648 = s_649 & s_662;
  assign s_649 = s_650[1];
  assign s_650 = {s_651,s_658};
  assign s_651 = s_652 & s_656;
  assign s_652 = ~s_653;
  assign s_653 = s_654[1];
  assign s_654 = s_655[3:2];
  assign s_655 = s_619[3:0];
  assign s_656 = ~s_657;
  assign s_657 = s_654[0];
  assign s_658 = s_659 & s_661;
  assign s_659 = ~s_660;
  assign s_660 = s_654[1];
  assign s_661 = s_654[0];
  assign s_662 = s_663[1];
  assign s_663 = {s_664,s_670};
  assign s_664 = s_665 & s_668;
  assign s_665 = ~s_666;
  assign s_666 = s_667[1];
  assign s_667 = s_655[1:0];
  assign s_668 = ~s_669;
  assign s_669 = s_667[0];
  assign s_670 = s_671 & s_673;
  assign s_671 = ~s_672;
  assign s_672 = s_667[1];
  assign s_673 = s_667[0];
  assign s_674 = {s_675,s_677};
  assign s_675 = s_649 & s_676;
  assign s_676 = ~s_662;
  assign s_677 = s_649?s_678:s_679;
  assign s_678 = s_663[0:0];
  assign s_679 = s_650[0:0];
  assign s_680 = {s_681,s_683};
  assign s_681 = s_609 & s_682;
  assign s_682 = ~s_646;
  assign s_683 = s_609?s_684:s_685;
  assign s_684 = s_647[1:0];
  assign s_685 = s_610[1:0];
  assign s_686 = s_687[3];
  assign s_687 = {s_688,s_758};
  assign s_688 = s_689 & s_724;
  assign s_689 = s_690[2];
  assign s_690 = {s_691,s_718};
  assign s_691 = s_692 & s_706;
  assign s_692 = s_693[1];
  assign s_693 = {s_694,s_702};
  assign s_694 = s_695 & s_700;
  assign s_695 = ~s_696;
  assign s_696 = s_697[1];
  assign s_697 = s_698[3:2];
  assign s_698 = s_699[7:4];
  assign s_699 = s_620[7:0];
  assign s_700 = ~s_701;
  assign s_701 = s_697[0];
  assign s_702 = s_703 & s_705;
  assign s_703 = ~s_704;
  assign s_704 = s_697[1];
  assign s_705 = s_697[0];
  assign s_706 = s_707[1];
  assign s_707 = {s_708,s_714};
  assign s_708 = s_709 & s_712;
  assign s_709 = ~s_710;
  assign s_710 = s_711[1];
  assign s_711 = s_698[1:0];
  assign s_712 = ~s_713;
  assign s_713 = s_711[0];
  assign s_714 = s_715 & s_717;
  assign s_715 = ~s_716;
  assign s_716 = s_711[1];
  assign s_717 = s_711[0];
  assign s_718 = {s_719,s_721};
  assign s_719 = s_692 & s_720;
  assign s_720 = ~s_706;
  assign s_721 = s_692?s_722:s_723;
  assign s_722 = s_707[0:0];
  assign s_723 = s_693[0:0];
  assign s_724 = s_725[2];
  assign s_725 = {s_726,s_752};
  assign s_726 = s_727 & s_740;
  assign s_727 = s_728[1];
  assign s_728 = {s_729,s_736};
  assign s_729 = s_730 & s_734;
  assign s_730 = ~s_731;
  assign s_731 = s_732[1];
  assign s_732 = s_733[3:2];
  assign s_733 = s_699[3:0];
  assign s_734 = ~s_735;
  assign s_735 = s_732[0];
  assign s_736 = s_737 & s_739;
  assign s_737 = ~s_738;
  assign s_738 = s_732[1];
  assign s_739 = s_732[0];
  assign s_740 = s_741[1];
  assign s_741 = {s_742,s_748};
  assign s_742 = s_743 & s_746;
  assign s_743 = ~s_744;
  assign s_744 = s_745[1];
  assign s_745 = s_733[1:0];
  assign s_746 = ~s_747;
  assign s_747 = s_745[0];
  assign s_748 = s_749 & s_751;
  assign s_749 = ~s_750;
  assign s_750 = s_745[1];
  assign s_751 = s_745[0];
  assign s_752 = {s_753,s_755};
  assign s_753 = s_727 & s_754;
  assign s_754 = ~s_740;
  assign s_755 = s_727?s_756:s_757;
  assign s_756 = s_741[0:0];
  assign s_757 = s_728[0:0];
  assign s_758 = {s_759,s_761};
  assign s_759 = s_689 & s_760;
  assign s_760 = ~s_724;
  assign s_761 = s_689?s_762:s_763;
  assign s_762 = s_725[1:0];
  assign s_763 = s_690[1:0];
  assign s_764 = {s_765,s_767};
  assign s_765 = s_606 & s_766;
  assign s_766 = ~s_686;
  assign s_767 = s_606?s_768:s_769;
  assign s_768 = s_687[2:0];
  assign s_769 = s_607[2:0];
  assign s_770 = s_771[4];
  assign s_771 = {s_772,s_930};
  assign s_772 = s_773 & s_852;
  assign s_773 = s_774[3];
  assign s_774 = {s_775,s_846};
  assign s_775 = s_776 & s_812;
  assign s_776 = s_777[2];
  assign s_777 = {s_778,s_806};
  assign s_778 = s_779 & s_794;
  assign s_779 = s_780[1];
  assign s_780 = {s_781,s_790};
  assign s_781 = s_782 & s_788;
  assign s_782 = ~s_783;
  assign s_783 = s_784[1];
  assign s_784 = s_785[3:2];
  assign s_785 = s_786[7:4];
  assign s_786 = s_787[15:8];
  assign s_787 = s_621[15:0];
  assign s_788 = ~s_789;
  assign s_789 = s_784[0];
  assign s_790 = s_791 & s_793;
  assign s_791 = ~s_792;
  assign s_792 = s_784[1];
  assign s_793 = s_784[0];
  assign s_794 = s_795[1];
  assign s_795 = {s_796,s_802};
  assign s_796 = s_797 & s_800;
  assign s_797 = ~s_798;
  assign s_798 = s_799[1];
  assign s_799 = s_785[1:0];
  assign s_800 = ~s_801;
  assign s_801 = s_799[0];
  assign s_802 = s_803 & s_805;
  assign s_803 = ~s_804;
  assign s_804 = s_799[1];
  assign s_805 = s_799[0];
  assign s_806 = {s_807,s_809};
  assign s_807 = s_779 & s_808;
  assign s_808 = ~s_794;
  assign s_809 = s_779?s_810:s_811;
  assign s_810 = s_795[0:0];
  assign s_811 = s_780[0:0];
  assign s_812 = s_813[2];
  assign s_813 = {s_814,s_840};
  assign s_814 = s_815 & s_828;
  assign s_815 = s_816[1];
  assign s_816 = {s_817,s_824};
  assign s_817 = s_818 & s_822;
  assign s_818 = ~s_819;
  assign s_819 = s_820[1];
  assign s_820 = s_821[3:2];
  assign s_821 = s_786[3:0];
  assign s_822 = ~s_823;
  assign s_823 = s_820[0];
  assign s_824 = s_825 & s_827;
  assign s_825 = ~s_826;
  assign s_826 = s_820[1];
  assign s_827 = s_820[0];
  assign s_828 = s_829[1];
  assign s_829 = {s_830,s_836};
  assign s_830 = s_831 & s_834;
  assign s_831 = ~s_832;
  assign s_832 = s_833[1];
  assign s_833 = s_821[1:0];
  assign s_834 = ~s_835;
  assign s_835 = s_833[0];
  assign s_836 = s_837 & s_839;
  assign s_837 = ~s_838;
  assign s_838 = s_833[1];
  assign s_839 = s_833[0];
  assign s_840 = {s_841,s_843};
  assign s_841 = s_815 & s_842;
  assign s_842 = ~s_828;
  assign s_843 = s_815?s_844:s_845;
  assign s_844 = s_829[0:0];
  assign s_845 = s_816[0:0];
  assign s_846 = {s_847,s_849};
  assign s_847 = s_776 & s_848;
  assign s_848 = ~s_812;
  assign s_849 = s_776?s_850:s_851;
  assign s_850 = s_813[1:0];
  assign s_851 = s_777[1:0];
  assign s_852 = s_853[3];
  assign s_853 = {s_854,s_924};
  assign s_854 = s_855 & s_890;
  assign s_855 = s_856[2];
  assign s_856 = {s_857,s_884};
  assign s_857 = s_858 & s_872;
  assign s_858 = s_859[1];
  assign s_859 = {s_860,s_868};
  assign s_860 = s_861 & s_866;
  assign s_861 = ~s_862;
  assign s_862 = s_863[1];
  assign s_863 = s_864[3:2];
  assign s_864 = s_865[7:4];
  assign s_865 = s_787[7:0];
  assign s_866 = ~s_867;
  assign s_867 = s_863[0];
  assign s_868 = s_869 & s_871;
  assign s_869 = ~s_870;
  assign s_870 = s_863[1];
  assign s_871 = s_863[0];
  assign s_872 = s_873[1];
  assign s_873 = {s_874,s_880};
  assign s_874 = s_875 & s_878;
  assign s_875 = ~s_876;
  assign s_876 = s_877[1];
  assign s_877 = s_864[1:0];
  assign s_878 = ~s_879;
  assign s_879 = s_877[0];
  assign s_880 = s_881 & s_883;
  assign s_881 = ~s_882;
  assign s_882 = s_877[1];
  assign s_883 = s_877[0];
  assign s_884 = {s_885,s_887};
  assign s_885 = s_858 & s_886;
  assign s_886 = ~s_872;
  assign s_887 = s_858?s_888:s_889;
  assign s_888 = s_873[0:0];
  assign s_889 = s_859[0:0];
  assign s_890 = s_891[2];
  assign s_891 = {s_892,s_918};
  assign s_892 = s_893 & s_906;
  assign s_893 = s_894[1];
  assign s_894 = {s_895,s_902};
  assign s_895 = s_896 & s_900;
  assign s_896 = ~s_897;
  assign s_897 = s_898[1];
  assign s_898 = s_899[3:2];
  assign s_899 = s_865[3:0];
  assign s_900 = ~s_901;
  assign s_901 = s_898[0];
  assign s_902 = s_903 & s_905;
  assign s_903 = ~s_904;
  assign s_904 = s_898[1];
  assign s_905 = s_898[0];
  assign s_906 = s_907[1];
  assign s_907 = {s_908,s_914};
  assign s_908 = s_909 & s_912;
  assign s_909 = ~s_910;
  assign s_910 = s_911[1];
  assign s_911 = s_899[1:0];
  assign s_912 = ~s_913;
  assign s_913 = s_911[0];
  assign s_914 = s_915 & s_917;
  assign s_915 = ~s_916;
  assign s_916 = s_911[1];
  assign s_917 = s_911[0];
  assign s_918 = {s_919,s_921};
  assign s_919 = s_893 & s_920;
  assign s_920 = ~s_906;
  assign s_921 = s_893?s_922:s_923;
  assign s_922 = s_907[0:0];
  assign s_923 = s_894[0:0];
  assign s_924 = {s_925,s_927};
  assign s_925 = s_855 & s_926;
  assign s_926 = ~s_890;
  assign s_927 = s_855?s_928:s_929;
  assign s_928 = s_891[1:0];
  assign s_929 = s_856[1:0];
  assign s_930 = {s_931,s_933};
  assign s_931 = s_773 & s_932;
  assign s_932 = ~s_852;
  assign s_933 = s_773?s_934:s_935;
  assign s_934 = s_853[2:0];
  assign s_935 = s_774[2:0];
  assign s_936 = {s_937,s_939};
  assign s_937 = s_603 & s_938;
  assign s_938 = ~s_770;
  assign s_939 = s_603?s_940:s_941;
  assign s_940 = s_771[3:0];
  assign s_941 = s_604[3:0];
  assign s_942 = {s_943,s_945};
  assign s_943 = s_236 & s_944;
  assign s_944 = ~s_600;
  assign s_945 = s_236?s_946:s_947;
  assign s_946 = s_601[4:0];
  assign s_947 = s_237[4:0];
  dq #(13, 1) dq_s_948 (clk, s_948, s_949);
  assign s_949 = s_950 - s_953;
  assign s_950 = $signed(s_951);
  assign s_951 = s_225?s_952:s_226;
  assign s_952 = -11'd1022;
  assign s_953 = -13'd2044;
  assign s_954 = s_955 <= s_956;
  assign s_955 = s_233;
  dq #(13, 1) dq_s_956 (clk, s_956, s_949);
  assign s_957 = 2'd3;
  assign s_958 = s_959 << s_1699;
  assign s_959 = s_960;
  dq #(53, 1) dq_s_960 (clk, s_960, s_961);
  assign s_961 = s_962 << s_973;
  dq #(53, 2) dq_s_962 (clk, s_962, s_963);
  assign s_963 = {s_964,s_972};
  assign s_964 = s_967?s_965:s_966;
  assign s_965 = 1'd0;
  assign s_966 = 1'd1;
  assign s_967 = s_968 == s_971;
  assign s_968 = s_969 - s_970;
  assign s_969 = s_7[62:52];
  assign s_970 = 10'd1023;
  assign s_971 = -11'd1023;
  assign s_972 = s_7[51:0];
  dq #(13, 1) dq_s_973 (clk, s_973, s_974);
  assign s_974 = s_1696?s_975:s_1690;
  dq #(7, 1) dq_s_975 (clk, s_975, s_976);
  assign s_976 = {s_977,s_1684};
  assign s_977 = s_978 & s_1342;
  assign s_978 = s_979[5];
  assign s_979 = {s_980,s_1336};
  assign s_980 = s_981 & s_1170;
  assign s_981 = s_982[4];
  assign s_982 = {s_983,s_1164};
  assign s_983 = s_984 & s_1086;
  assign s_984 = s_985[3];
  assign s_985 = {s_986,s_1080};
  assign s_986 = s_987 & s_1046;
  assign s_987 = s_988[2];
  assign s_988 = {s_989,s_1040};
  assign s_989 = s_990 & s_1028;
  assign s_990 = s_991[1];
  assign s_991 = {s_992,s_1024};
  assign s_992 = s_993 & s_1022;
  assign s_993 = ~s_994;
  assign s_994 = s_995[1];
  assign s_995 = s_996[3:2];
  assign s_996 = s_997[7:4];
  assign s_997 = s_998[15:8];
  assign s_998 = s_999[31:16];
  assign s_999 = s_1000[63:32];
  assign s_1000 = {s_1001,s_1021};
  assign s_1001 = {s_1002,s_1020};
  assign s_1002 = {s_1003,s_1019};
  assign s_1003 = {s_1004,s_1018};
  assign s_1004 = {s_1005,s_1017};
  assign s_1005 = {s_1006,s_1016};
  assign s_1006 = {s_1007,s_1015};
  assign s_1007 = {s_1008,s_1014};
  assign s_1008 = {s_1009,s_1013};
  assign s_1009 = {s_1010,s_1012};
  assign s_1010 = {s_963,s_1011};
  assign s_1011 = 1'd1;
  assign s_1012 = 1'd1;
  assign s_1013 = 1'd1;
  assign s_1014 = 1'd1;
  assign s_1015 = 1'd1;
  assign s_1016 = 1'd1;
  assign s_1017 = 1'd1;
  assign s_1018 = 1'd1;
  assign s_1019 = 1'd1;
  assign s_1020 = 1'd1;
  assign s_1021 = 1'd1;
  assign s_1022 = ~s_1023;
  assign s_1023 = s_995[0];
  assign s_1024 = s_1025 & s_1027;
  assign s_1025 = ~s_1026;
  assign s_1026 = s_995[1];
  assign s_1027 = s_995[0];
  assign s_1028 = s_1029[1];
  assign s_1029 = {s_1030,s_1036};
  assign s_1030 = s_1031 & s_1034;
  assign s_1031 = ~s_1032;
  assign s_1032 = s_1033[1];
  assign s_1033 = s_996[1:0];
  assign s_1034 = ~s_1035;
  assign s_1035 = s_1033[0];
  assign s_1036 = s_1037 & s_1039;
  assign s_1037 = ~s_1038;
  assign s_1038 = s_1033[1];
  assign s_1039 = s_1033[0];
  assign s_1040 = {s_1041,s_1043};
  assign s_1041 = s_990 & s_1042;
  assign s_1042 = ~s_1028;
  assign s_1043 = s_990?s_1044:s_1045;
  assign s_1044 = s_1029[0:0];
  assign s_1045 = s_991[0:0];
  assign s_1046 = s_1047[2];
  assign s_1047 = {s_1048,s_1074};
  assign s_1048 = s_1049 & s_1062;
  assign s_1049 = s_1050[1];
  assign s_1050 = {s_1051,s_1058};
  assign s_1051 = s_1052 & s_1056;
  assign s_1052 = ~s_1053;
  assign s_1053 = s_1054[1];
  assign s_1054 = s_1055[3:2];
  assign s_1055 = s_997[3:0];
  assign s_1056 = ~s_1057;
  assign s_1057 = s_1054[0];
  assign s_1058 = s_1059 & s_1061;
  assign s_1059 = ~s_1060;
  assign s_1060 = s_1054[1];
  assign s_1061 = s_1054[0];
  assign s_1062 = s_1063[1];
  assign s_1063 = {s_1064,s_1070};
  assign s_1064 = s_1065 & s_1068;
  assign s_1065 = ~s_1066;
  assign s_1066 = s_1067[1];
  assign s_1067 = s_1055[1:0];
  assign s_1068 = ~s_1069;
  assign s_1069 = s_1067[0];
  assign s_1070 = s_1071 & s_1073;
  assign s_1071 = ~s_1072;
  assign s_1072 = s_1067[1];
  assign s_1073 = s_1067[0];
  assign s_1074 = {s_1075,s_1077};
  assign s_1075 = s_1049 & s_1076;
  assign s_1076 = ~s_1062;
  assign s_1077 = s_1049?s_1078:s_1079;
  assign s_1078 = s_1063[0:0];
  assign s_1079 = s_1050[0:0];
  assign s_1080 = {s_1081,s_1083};
  assign s_1081 = s_987 & s_1082;
  assign s_1082 = ~s_1046;
  assign s_1083 = s_987?s_1084:s_1085;
  assign s_1084 = s_1047[1:0];
  assign s_1085 = s_988[1:0];
  assign s_1086 = s_1087[3];
  assign s_1087 = {s_1088,s_1158};
  assign s_1088 = s_1089 & s_1124;
  assign s_1089 = s_1090[2];
  assign s_1090 = {s_1091,s_1118};
  assign s_1091 = s_1092 & s_1106;
  assign s_1092 = s_1093[1];
  assign s_1093 = {s_1094,s_1102};
  assign s_1094 = s_1095 & s_1100;
  assign s_1095 = ~s_1096;
  assign s_1096 = s_1097[1];
  assign s_1097 = s_1098[3:2];
  assign s_1098 = s_1099[7:4];
  assign s_1099 = s_998[7:0];
  assign s_1100 = ~s_1101;
  assign s_1101 = s_1097[0];
  assign s_1102 = s_1103 & s_1105;
  assign s_1103 = ~s_1104;
  assign s_1104 = s_1097[1];
  assign s_1105 = s_1097[0];
  assign s_1106 = s_1107[1];
  assign s_1107 = {s_1108,s_1114};
  assign s_1108 = s_1109 & s_1112;
  assign s_1109 = ~s_1110;
  assign s_1110 = s_1111[1];
  assign s_1111 = s_1098[1:0];
  assign s_1112 = ~s_1113;
  assign s_1113 = s_1111[0];
  assign s_1114 = s_1115 & s_1117;
  assign s_1115 = ~s_1116;
  assign s_1116 = s_1111[1];
  assign s_1117 = s_1111[0];
  assign s_1118 = {s_1119,s_1121};
  assign s_1119 = s_1092 & s_1120;
  assign s_1120 = ~s_1106;
  assign s_1121 = s_1092?s_1122:s_1123;
  assign s_1122 = s_1107[0:0];
  assign s_1123 = s_1093[0:0];
  assign s_1124 = s_1125[2];
  assign s_1125 = {s_1126,s_1152};
  assign s_1126 = s_1127 & s_1140;
  assign s_1127 = s_1128[1];
  assign s_1128 = {s_1129,s_1136};
  assign s_1129 = s_1130 & s_1134;
  assign s_1130 = ~s_1131;
  assign s_1131 = s_1132[1];
  assign s_1132 = s_1133[3:2];
  assign s_1133 = s_1099[3:0];
  assign s_1134 = ~s_1135;
  assign s_1135 = s_1132[0];
  assign s_1136 = s_1137 & s_1139;
  assign s_1137 = ~s_1138;
  assign s_1138 = s_1132[1];
  assign s_1139 = s_1132[0];
  assign s_1140 = s_1141[1];
  assign s_1141 = {s_1142,s_1148};
  assign s_1142 = s_1143 & s_1146;
  assign s_1143 = ~s_1144;
  assign s_1144 = s_1145[1];
  assign s_1145 = s_1133[1:0];
  assign s_1146 = ~s_1147;
  assign s_1147 = s_1145[0];
  assign s_1148 = s_1149 & s_1151;
  assign s_1149 = ~s_1150;
  assign s_1150 = s_1145[1];
  assign s_1151 = s_1145[0];
  assign s_1152 = {s_1153,s_1155};
  assign s_1153 = s_1127 & s_1154;
  assign s_1154 = ~s_1140;
  assign s_1155 = s_1127?s_1156:s_1157;
  assign s_1156 = s_1141[0:0];
  assign s_1157 = s_1128[0:0];
  assign s_1158 = {s_1159,s_1161};
  assign s_1159 = s_1089 & s_1160;
  assign s_1160 = ~s_1124;
  assign s_1161 = s_1089?s_1162:s_1163;
  assign s_1162 = s_1125[1:0];
  assign s_1163 = s_1090[1:0];
  assign s_1164 = {s_1165,s_1167};
  assign s_1165 = s_984 & s_1166;
  assign s_1166 = ~s_1086;
  assign s_1167 = s_984?s_1168:s_1169;
  assign s_1168 = s_1087[2:0];
  assign s_1169 = s_985[2:0];
  assign s_1170 = s_1171[4];
  assign s_1171 = {s_1172,s_1330};
  assign s_1172 = s_1173 & s_1252;
  assign s_1173 = s_1174[3];
  assign s_1174 = {s_1175,s_1246};
  assign s_1175 = s_1176 & s_1212;
  assign s_1176 = s_1177[2];
  assign s_1177 = {s_1178,s_1206};
  assign s_1178 = s_1179 & s_1194;
  assign s_1179 = s_1180[1];
  assign s_1180 = {s_1181,s_1190};
  assign s_1181 = s_1182 & s_1188;
  assign s_1182 = ~s_1183;
  assign s_1183 = s_1184[1];
  assign s_1184 = s_1185[3:2];
  assign s_1185 = s_1186[7:4];
  assign s_1186 = s_1187[15:8];
  assign s_1187 = s_999[15:0];
  assign s_1188 = ~s_1189;
  assign s_1189 = s_1184[0];
  assign s_1190 = s_1191 & s_1193;
  assign s_1191 = ~s_1192;
  assign s_1192 = s_1184[1];
  assign s_1193 = s_1184[0];
  assign s_1194 = s_1195[1];
  assign s_1195 = {s_1196,s_1202};
  assign s_1196 = s_1197 & s_1200;
  assign s_1197 = ~s_1198;
  assign s_1198 = s_1199[1];
  assign s_1199 = s_1185[1:0];
  assign s_1200 = ~s_1201;
  assign s_1201 = s_1199[0];
  assign s_1202 = s_1203 & s_1205;
  assign s_1203 = ~s_1204;
  assign s_1204 = s_1199[1];
  assign s_1205 = s_1199[0];
  assign s_1206 = {s_1207,s_1209};
  assign s_1207 = s_1179 & s_1208;
  assign s_1208 = ~s_1194;
  assign s_1209 = s_1179?s_1210:s_1211;
  assign s_1210 = s_1195[0:0];
  assign s_1211 = s_1180[0:0];
  assign s_1212 = s_1213[2];
  assign s_1213 = {s_1214,s_1240};
  assign s_1214 = s_1215 & s_1228;
  assign s_1215 = s_1216[1];
  assign s_1216 = {s_1217,s_1224};
  assign s_1217 = s_1218 & s_1222;
  assign s_1218 = ~s_1219;
  assign s_1219 = s_1220[1];
  assign s_1220 = s_1221[3:2];
  assign s_1221 = s_1186[3:0];
  assign s_1222 = ~s_1223;
  assign s_1223 = s_1220[0];
  assign s_1224 = s_1225 & s_1227;
  assign s_1225 = ~s_1226;
  assign s_1226 = s_1220[1];
  assign s_1227 = s_1220[0];
  assign s_1228 = s_1229[1];
  assign s_1229 = {s_1230,s_1236};
  assign s_1230 = s_1231 & s_1234;
  assign s_1231 = ~s_1232;
  assign s_1232 = s_1233[1];
  assign s_1233 = s_1221[1:0];
  assign s_1234 = ~s_1235;
  assign s_1235 = s_1233[0];
  assign s_1236 = s_1237 & s_1239;
  assign s_1237 = ~s_1238;
  assign s_1238 = s_1233[1];
  assign s_1239 = s_1233[0];
  assign s_1240 = {s_1241,s_1243};
  assign s_1241 = s_1215 & s_1242;
  assign s_1242 = ~s_1228;
  assign s_1243 = s_1215?s_1244:s_1245;
  assign s_1244 = s_1229[0:0];
  assign s_1245 = s_1216[0:0];
  assign s_1246 = {s_1247,s_1249};
  assign s_1247 = s_1176 & s_1248;
  assign s_1248 = ~s_1212;
  assign s_1249 = s_1176?s_1250:s_1251;
  assign s_1250 = s_1213[1:0];
  assign s_1251 = s_1177[1:0];
  assign s_1252 = s_1253[3];
  assign s_1253 = {s_1254,s_1324};
  assign s_1254 = s_1255 & s_1290;
  assign s_1255 = s_1256[2];
  assign s_1256 = {s_1257,s_1284};
  assign s_1257 = s_1258 & s_1272;
  assign s_1258 = s_1259[1];
  assign s_1259 = {s_1260,s_1268};
  assign s_1260 = s_1261 & s_1266;
  assign s_1261 = ~s_1262;
  assign s_1262 = s_1263[1];
  assign s_1263 = s_1264[3:2];
  assign s_1264 = s_1265[7:4];
  assign s_1265 = s_1187[7:0];
  assign s_1266 = ~s_1267;
  assign s_1267 = s_1263[0];
  assign s_1268 = s_1269 & s_1271;
  assign s_1269 = ~s_1270;
  assign s_1270 = s_1263[1];
  assign s_1271 = s_1263[0];
  assign s_1272 = s_1273[1];
  assign s_1273 = {s_1274,s_1280};
  assign s_1274 = s_1275 & s_1278;
  assign s_1275 = ~s_1276;
  assign s_1276 = s_1277[1];
  assign s_1277 = s_1264[1:0];
  assign s_1278 = ~s_1279;
  assign s_1279 = s_1277[0];
  assign s_1280 = s_1281 & s_1283;
  assign s_1281 = ~s_1282;
  assign s_1282 = s_1277[1];
  assign s_1283 = s_1277[0];
  assign s_1284 = {s_1285,s_1287};
  assign s_1285 = s_1258 & s_1286;
  assign s_1286 = ~s_1272;
  assign s_1287 = s_1258?s_1288:s_1289;
  assign s_1288 = s_1273[0:0];
  assign s_1289 = s_1259[0:0];
  assign s_1290 = s_1291[2];
  assign s_1291 = {s_1292,s_1318};
  assign s_1292 = s_1293 & s_1306;
  assign s_1293 = s_1294[1];
  assign s_1294 = {s_1295,s_1302};
  assign s_1295 = s_1296 & s_1300;
  assign s_1296 = ~s_1297;
  assign s_1297 = s_1298[1];
  assign s_1298 = s_1299[3:2];
  assign s_1299 = s_1265[3:0];
  assign s_1300 = ~s_1301;
  assign s_1301 = s_1298[0];
  assign s_1302 = s_1303 & s_1305;
  assign s_1303 = ~s_1304;
  assign s_1304 = s_1298[1];
  assign s_1305 = s_1298[0];
  assign s_1306 = s_1307[1];
  assign s_1307 = {s_1308,s_1314};
  assign s_1308 = s_1309 & s_1312;
  assign s_1309 = ~s_1310;
  assign s_1310 = s_1311[1];
  assign s_1311 = s_1299[1:0];
  assign s_1312 = ~s_1313;
  assign s_1313 = s_1311[0];
  assign s_1314 = s_1315 & s_1317;
  assign s_1315 = ~s_1316;
  assign s_1316 = s_1311[1];
  assign s_1317 = s_1311[0];
  assign s_1318 = {s_1319,s_1321};
  assign s_1319 = s_1293 & s_1320;
  assign s_1320 = ~s_1306;
  assign s_1321 = s_1293?s_1322:s_1323;
  assign s_1322 = s_1307[0:0];
  assign s_1323 = s_1294[0:0];
  assign s_1324 = {s_1325,s_1327};
  assign s_1325 = s_1255 & s_1326;
  assign s_1326 = ~s_1290;
  assign s_1327 = s_1255?s_1328:s_1329;
  assign s_1328 = s_1291[1:0];
  assign s_1329 = s_1256[1:0];
  assign s_1330 = {s_1331,s_1333};
  assign s_1331 = s_1173 & s_1332;
  assign s_1332 = ~s_1252;
  assign s_1333 = s_1173?s_1334:s_1335;
  assign s_1334 = s_1253[2:0];
  assign s_1335 = s_1174[2:0];
  assign s_1336 = {s_1337,s_1339};
  assign s_1337 = s_981 & s_1338;
  assign s_1338 = ~s_1170;
  assign s_1339 = s_981?s_1340:s_1341;
  assign s_1340 = s_1171[3:0];
  assign s_1341 = s_982[3:0];
  assign s_1342 = s_1343[5];
  assign s_1343 = {s_1344,s_1678};
  assign s_1344 = s_1345 & s_1512;
  assign s_1345 = s_1346[4];
  assign s_1346 = {s_1347,s_1506};
  assign s_1347 = s_1348 & s_1428;
  assign s_1348 = s_1349[3];
  assign s_1349 = {s_1350,s_1422};
  assign s_1350 = s_1351 & s_1388;
  assign s_1351 = s_1352[2];
  assign s_1352 = {s_1353,s_1382};
  assign s_1353 = s_1354 & s_1370;
  assign s_1354 = s_1355[1];
  assign s_1355 = {s_1356,s_1366};
  assign s_1356 = s_1357 & s_1364;
  assign s_1357 = ~s_1358;
  assign s_1358 = s_1359[1];
  assign s_1359 = s_1360[3:2];
  assign s_1360 = s_1361[7:4];
  assign s_1361 = s_1362[15:8];
  assign s_1362 = s_1363[31:16];
  assign s_1363 = s_1000[31:0];
  assign s_1364 = ~s_1365;
  assign s_1365 = s_1359[0];
  assign s_1366 = s_1367 & s_1369;
  assign s_1367 = ~s_1368;
  assign s_1368 = s_1359[1];
  assign s_1369 = s_1359[0];
  assign s_1370 = s_1371[1];
  assign s_1371 = {s_1372,s_1378};
  assign s_1372 = s_1373 & s_1376;
  assign s_1373 = ~s_1374;
  assign s_1374 = s_1375[1];
  assign s_1375 = s_1360[1:0];
  assign s_1376 = ~s_1377;
  assign s_1377 = s_1375[0];
  assign s_1378 = s_1379 & s_1381;
  assign s_1379 = ~s_1380;
  assign s_1380 = s_1375[1];
  assign s_1381 = s_1375[0];
  assign s_1382 = {s_1383,s_1385};
  assign s_1383 = s_1354 & s_1384;
  assign s_1384 = ~s_1370;
  assign s_1385 = s_1354?s_1386:s_1387;
  assign s_1386 = s_1371[0:0];
  assign s_1387 = s_1355[0:0];
  assign s_1388 = s_1389[2];
  assign s_1389 = {s_1390,s_1416};
  assign s_1390 = s_1391 & s_1404;
  assign s_1391 = s_1392[1];
  assign s_1392 = {s_1393,s_1400};
  assign s_1393 = s_1394 & s_1398;
  assign s_1394 = ~s_1395;
  assign s_1395 = s_1396[1];
  assign s_1396 = s_1397[3:2];
  assign s_1397 = s_1361[3:0];
  assign s_1398 = ~s_1399;
  assign s_1399 = s_1396[0];
  assign s_1400 = s_1401 & s_1403;
  assign s_1401 = ~s_1402;
  assign s_1402 = s_1396[1];
  assign s_1403 = s_1396[0];
  assign s_1404 = s_1405[1];
  assign s_1405 = {s_1406,s_1412};
  assign s_1406 = s_1407 & s_1410;
  assign s_1407 = ~s_1408;
  assign s_1408 = s_1409[1];
  assign s_1409 = s_1397[1:0];
  assign s_1410 = ~s_1411;
  assign s_1411 = s_1409[0];
  assign s_1412 = s_1413 & s_1415;
  assign s_1413 = ~s_1414;
  assign s_1414 = s_1409[1];
  assign s_1415 = s_1409[0];
  assign s_1416 = {s_1417,s_1419};
  assign s_1417 = s_1391 & s_1418;
  assign s_1418 = ~s_1404;
  assign s_1419 = s_1391?s_1420:s_1421;
  assign s_1420 = s_1405[0:0];
  assign s_1421 = s_1392[0:0];
  assign s_1422 = {s_1423,s_1425};
  assign s_1423 = s_1351 & s_1424;
  assign s_1424 = ~s_1388;
  assign s_1425 = s_1351?s_1426:s_1427;
  assign s_1426 = s_1389[1:0];
  assign s_1427 = s_1352[1:0];
  assign s_1428 = s_1429[3];
  assign s_1429 = {s_1430,s_1500};
  assign s_1430 = s_1431 & s_1466;
  assign s_1431 = s_1432[2];
  assign s_1432 = {s_1433,s_1460};
  assign s_1433 = s_1434 & s_1448;
  assign s_1434 = s_1435[1];
  assign s_1435 = {s_1436,s_1444};
  assign s_1436 = s_1437 & s_1442;
  assign s_1437 = ~s_1438;
  assign s_1438 = s_1439[1];
  assign s_1439 = s_1440[3:2];
  assign s_1440 = s_1441[7:4];
  assign s_1441 = s_1362[7:0];
  assign s_1442 = ~s_1443;
  assign s_1443 = s_1439[0];
  assign s_1444 = s_1445 & s_1447;
  assign s_1445 = ~s_1446;
  assign s_1446 = s_1439[1];
  assign s_1447 = s_1439[0];
  assign s_1448 = s_1449[1];
  assign s_1449 = {s_1450,s_1456};
  assign s_1450 = s_1451 & s_1454;
  assign s_1451 = ~s_1452;
  assign s_1452 = s_1453[1];
  assign s_1453 = s_1440[1:0];
  assign s_1454 = ~s_1455;
  assign s_1455 = s_1453[0];
  assign s_1456 = s_1457 & s_1459;
  assign s_1457 = ~s_1458;
  assign s_1458 = s_1453[1];
  assign s_1459 = s_1453[0];
  assign s_1460 = {s_1461,s_1463};
  assign s_1461 = s_1434 & s_1462;
  assign s_1462 = ~s_1448;
  assign s_1463 = s_1434?s_1464:s_1465;
  assign s_1464 = s_1449[0:0];
  assign s_1465 = s_1435[0:0];
  assign s_1466 = s_1467[2];
  assign s_1467 = {s_1468,s_1494};
  assign s_1468 = s_1469 & s_1482;
  assign s_1469 = s_1470[1];
  assign s_1470 = {s_1471,s_1478};
  assign s_1471 = s_1472 & s_1476;
  assign s_1472 = ~s_1473;
  assign s_1473 = s_1474[1];
  assign s_1474 = s_1475[3:2];
  assign s_1475 = s_1441[3:0];
  assign s_1476 = ~s_1477;
  assign s_1477 = s_1474[0];
  assign s_1478 = s_1479 & s_1481;
  assign s_1479 = ~s_1480;
  assign s_1480 = s_1474[1];
  assign s_1481 = s_1474[0];
  assign s_1482 = s_1483[1];
  assign s_1483 = {s_1484,s_1490};
  assign s_1484 = s_1485 & s_1488;
  assign s_1485 = ~s_1486;
  assign s_1486 = s_1487[1];
  assign s_1487 = s_1475[1:0];
  assign s_1488 = ~s_1489;
  assign s_1489 = s_1487[0];
  assign s_1490 = s_1491 & s_1493;
  assign s_1491 = ~s_1492;
  assign s_1492 = s_1487[1];
  assign s_1493 = s_1487[0];
  assign s_1494 = {s_1495,s_1497};
  assign s_1495 = s_1469 & s_1496;
  assign s_1496 = ~s_1482;
  assign s_1497 = s_1469?s_1498:s_1499;
  assign s_1498 = s_1483[0:0];
  assign s_1499 = s_1470[0:0];
  assign s_1500 = {s_1501,s_1503};
  assign s_1501 = s_1431 & s_1502;
  assign s_1502 = ~s_1466;
  assign s_1503 = s_1431?s_1504:s_1505;
  assign s_1504 = s_1467[1:0];
  assign s_1505 = s_1432[1:0];
  assign s_1506 = {s_1507,s_1509};
  assign s_1507 = s_1348 & s_1508;
  assign s_1508 = ~s_1428;
  assign s_1509 = s_1348?s_1510:s_1511;
  assign s_1510 = s_1429[2:0];
  assign s_1511 = s_1349[2:0];
  assign s_1512 = s_1513[4];
  assign s_1513 = {s_1514,s_1672};
  assign s_1514 = s_1515 & s_1594;
  assign s_1515 = s_1516[3];
  assign s_1516 = {s_1517,s_1588};
  assign s_1517 = s_1518 & s_1554;
  assign s_1518 = s_1519[2];
  assign s_1519 = {s_1520,s_1548};
  assign s_1520 = s_1521 & s_1536;
  assign s_1521 = s_1522[1];
  assign s_1522 = {s_1523,s_1532};
  assign s_1523 = s_1524 & s_1530;
  assign s_1524 = ~s_1525;
  assign s_1525 = s_1526[1];
  assign s_1526 = s_1527[3:2];
  assign s_1527 = s_1528[7:4];
  assign s_1528 = s_1529[15:8];
  assign s_1529 = s_1363[15:0];
  assign s_1530 = ~s_1531;
  assign s_1531 = s_1526[0];
  assign s_1532 = s_1533 & s_1535;
  assign s_1533 = ~s_1534;
  assign s_1534 = s_1526[1];
  assign s_1535 = s_1526[0];
  assign s_1536 = s_1537[1];
  assign s_1537 = {s_1538,s_1544};
  assign s_1538 = s_1539 & s_1542;
  assign s_1539 = ~s_1540;
  assign s_1540 = s_1541[1];
  assign s_1541 = s_1527[1:0];
  assign s_1542 = ~s_1543;
  assign s_1543 = s_1541[0];
  assign s_1544 = s_1545 & s_1547;
  assign s_1545 = ~s_1546;
  assign s_1546 = s_1541[1];
  assign s_1547 = s_1541[0];
  assign s_1548 = {s_1549,s_1551};
  assign s_1549 = s_1521 & s_1550;
  assign s_1550 = ~s_1536;
  assign s_1551 = s_1521?s_1552:s_1553;
  assign s_1552 = s_1537[0:0];
  assign s_1553 = s_1522[0:0];
  assign s_1554 = s_1555[2];
  assign s_1555 = {s_1556,s_1582};
  assign s_1556 = s_1557 & s_1570;
  assign s_1557 = s_1558[1];
  assign s_1558 = {s_1559,s_1566};
  assign s_1559 = s_1560 & s_1564;
  assign s_1560 = ~s_1561;
  assign s_1561 = s_1562[1];
  assign s_1562 = s_1563[3:2];
  assign s_1563 = s_1528[3:0];
  assign s_1564 = ~s_1565;
  assign s_1565 = s_1562[0];
  assign s_1566 = s_1567 & s_1569;
  assign s_1567 = ~s_1568;
  assign s_1568 = s_1562[1];
  assign s_1569 = s_1562[0];
  assign s_1570 = s_1571[1];
  assign s_1571 = {s_1572,s_1578};
  assign s_1572 = s_1573 & s_1576;
  assign s_1573 = ~s_1574;
  assign s_1574 = s_1575[1];
  assign s_1575 = s_1563[1:0];
  assign s_1576 = ~s_1577;
  assign s_1577 = s_1575[0];
  assign s_1578 = s_1579 & s_1581;
  assign s_1579 = ~s_1580;
  assign s_1580 = s_1575[1];
  assign s_1581 = s_1575[0];
  assign s_1582 = {s_1583,s_1585};
  assign s_1583 = s_1557 & s_1584;
  assign s_1584 = ~s_1570;
  assign s_1585 = s_1557?s_1586:s_1587;
  assign s_1586 = s_1571[0:0];
  assign s_1587 = s_1558[0:0];
  assign s_1588 = {s_1589,s_1591};
  assign s_1589 = s_1518 & s_1590;
  assign s_1590 = ~s_1554;
  assign s_1591 = s_1518?s_1592:s_1593;
  assign s_1592 = s_1555[1:0];
  assign s_1593 = s_1519[1:0];
  assign s_1594 = s_1595[3];
  assign s_1595 = {s_1596,s_1666};
  assign s_1596 = s_1597 & s_1632;
  assign s_1597 = s_1598[2];
  assign s_1598 = {s_1599,s_1626};
  assign s_1599 = s_1600 & s_1614;
  assign s_1600 = s_1601[1];
  assign s_1601 = {s_1602,s_1610};
  assign s_1602 = s_1603 & s_1608;
  assign s_1603 = ~s_1604;
  assign s_1604 = s_1605[1];
  assign s_1605 = s_1606[3:2];
  assign s_1606 = s_1607[7:4];
  assign s_1607 = s_1529[7:0];
  assign s_1608 = ~s_1609;
  assign s_1609 = s_1605[0];
  assign s_1610 = s_1611 & s_1613;
  assign s_1611 = ~s_1612;
  assign s_1612 = s_1605[1];
  assign s_1613 = s_1605[0];
  assign s_1614 = s_1615[1];
  assign s_1615 = {s_1616,s_1622};
  assign s_1616 = s_1617 & s_1620;
  assign s_1617 = ~s_1618;
  assign s_1618 = s_1619[1];
  assign s_1619 = s_1606[1:0];
  assign s_1620 = ~s_1621;
  assign s_1621 = s_1619[0];
  assign s_1622 = s_1623 & s_1625;
  assign s_1623 = ~s_1624;
  assign s_1624 = s_1619[1];
  assign s_1625 = s_1619[0];
  assign s_1626 = {s_1627,s_1629};
  assign s_1627 = s_1600 & s_1628;
  assign s_1628 = ~s_1614;
  assign s_1629 = s_1600?s_1630:s_1631;
  assign s_1630 = s_1615[0:0];
  assign s_1631 = s_1601[0:0];
  assign s_1632 = s_1633[2];
  assign s_1633 = {s_1634,s_1660};
  assign s_1634 = s_1635 & s_1648;
  assign s_1635 = s_1636[1];
  assign s_1636 = {s_1637,s_1644};
  assign s_1637 = s_1638 & s_1642;
  assign s_1638 = ~s_1639;
  assign s_1639 = s_1640[1];
  assign s_1640 = s_1641[3:2];
  assign s_1641 = s_1607[3:0];
  assign s_1642 = ~s_1643;
  assign s_1643 = s_1640[0];
  assign s_1644 = s_1645 & s_1647;
  assign s_1645 = ~s_1646;
  assign s_1646 = s_1640[1];
  assign s_1647 = s_1640[0];
  assign s_1648 = s_1649[1];
  assign s_1649 = {s_1650,s_1656};
  assign s_1650 = s_1651 & s_1654;
  assign s_1651 = ~s_1652;
  assign s_1652 = s_1653[1];
  assign s_1653 = s_1641[1:0];
  assign s_1654 = ~s_1655;
  assign s_1655 = s_1653[0];
  assign s_1656 = s_1657 & s_1659;
  assign s_1657 = ~s_1658;
  assign s_1658 = s_1653[1];
  assign s_1659 = s_1653[0];
  assign s_1660 = {s_1661,s_1663};
  assign s_1661 = s_1635 & s_1662;
  assign s_1662 = ~s_1648;
  assign s_1663 = s_1635?s_1664:s_1665;
  assign s_1664 = s_1649[0:0];
  assign s_1665 = s_1636[0:0];
  assign s_1666 = {s_1667,s_1669};
  assign s_1667 = s_1597 & s_1668;
  assign s_1668 = ~s_1632;
  assign s_1669 = s_1597?s_1670:s_1671;
  assign s_1670 = s_1633[1:0];
  assign s_1671 = s_1598[1:0];
  assign s_1672 = {s_1673,s_1675};
  assign s_1673 = s_1515 & s_1674;
  assign s_1674 = ~s_1594;
  assign s_1675 = s_1515?s_1676:s_1677;
  assign s_1676 = s_1595[2:0];
  assign s_1677 = s_1516[2:0];
  assign s_1678 = {s_1679,s_1681};
  assign s_1679 = s_1345 & s_1680;
  assign s_1680 = ~s_1512;
  assign s_1681 = s_1345?s_1682:s_1683;
  assign s_1682 = s_1513[3:0];
  assign s_1683 = s_1346[3:0];
  assign s_1684 = {s_1685,s_1687};
  assign s_1685 = s_978 & s_1686;
  assign s_1686 = ~s_1342;
  assign s_1687 = s_978?s_1688:s_1689;
  assign s_1688 = s_1343[4:0];
  assign s_1689 = s_979[4:0];
  dq #(13, 1) dq_s_1690 (clk, s_1690, s_1691);
  assign s_1691 = s_1692 - s_1695;
  assign s_1692 = $signed(s_1693);
  assign s_1693 = s_967?s_1694:s_968;
  assign s_1694 = -11'd1022;
  assign s_1695 = -13'd2044;
  assign s_1696 = s_1697 <= s_1698;
  assign s_1697 = s_975;
  dq #(13, 1) dq_s_1698 (clk, s_1698, s_1691);
  assign s_1699 = 2'd3;
  assign s_1700 = 1'd1;
  assign s_1701 = s_203 | s_1702;
  assign s_1702 = 1'd1;
  assign s_1703 = s_1704[56];
  assign s_1704 = s_1705 - s_1712;
  assign s_1705 = s_1706;
  assign s_1706 = s_1707 | s_1711;
  assign s_1707 = s_1708 << s_1710;
  dq #(57, 1) dq_s_1708 (clk, s_1708, s_1709);
  assign s_1709 = s_213?s_216:s_214;
  assign s_1710 = 1'd1;
  assign s_1711 = 1'd0;
  dq #(56, 1) dq_s_1712 (clk, s_1712, s_958);
  assign s_1713 = 1'd1;
  assign s_1714 = s_200 | s_1715;
  assign s_1715 = 1'd1;
  assign s_1716 = s_1717[56];
  assign s_1717 = s_1718 - s_1725;
  assign s_1718 = s_1719;
  assign s_1719 = s_1720 | s_1724;
  assign s_1720 = s_1721 << s_1723;
  dq #(57, 1) dq_s_1721 (clk, s_1721, s_1722);
  assign s_1722 = s_1703?s_1706:s_1704;
  assign s_1723 = 1'd1;
  assign s_1724 = 1'd0;
  dq #(56, 2) dq_s_1725 (clk, s_1725, s_958);
  assign s_1726 = 1'd1;
  assign s_1727 = s_197 | s_1728;
  assign s_1728 = 1'd1;
  assign s_1729 = s_1730[56];
  assign s_1730 = s_1731 - s_1738;
  assign s_1731 = s_1732;
  assign s_1732 = s_1733 | s_1737;
  assign s_1733 = s_1734 << s_1736;
  dq #(57, 1) dq_s_1734 (clk, s_1734, s_1735);
  assign s_1735 = s_1716?s_1719:s_1717;
  assign s_1736 = 1'd1;
  assign s_1737 = 1'd0;
  dq #(56, 3) dq_s_1738 (clk, s_1738, s_958);
  assign s_1739 = 1'd1;
  assign s_1740 = s_194 | s_1741;
  assign s_1741 = 1'd1;
  assign s_1742 = s_1743[56];
  assign s_1743 = s_1744 - s_1751;
  assign s_1744 = s_1745;
  assign s_1745 = s_1746 | s_1750;
  assign s_1746 = s_1747 << s_1749;
  dq #(57, 1) dq_s_1747 (clk, s_1747, s_1748);
  assign s_1748 = s_1729?s_1732:s_1730;
  assign s_1749 = 1'd1;
  assign s_1750 = 1'd0;
  dq #(56, 4) dq_s_1751 (clk, s_1751, s_958);
  assign s_1752 = 1'd1;
  assign s_1753 = s_191 | s_1754;
  assign s_1754 = 1'd1;
  assign s_1755 = s_1756[56];
  assign s_1756 = s_1757 - s_1764;
  assign s_1757 = s_1758;
  assign s_1758 = s_1759 | s_1763;
  assign s_1759 = s_1760 << s_1762;
  dq #(57, 1) dq_s_1760 (clk, s_1760, s_1761);
  assign s_1761 = s_1742?s_1745:s_1743;
  assign s_1762 = 1'd1;
  assign s_1763 = 1'd0;
  dq #(56, 5) dq_s_1764 (clk, s_1764, s_958);
  assign s_1765 = 1'd1;
  assign s_1766 = s_188 | s_1767;
  assign s_1767 = 1'd1;
  assign s_1768 = s_1769[56];
  assign s_1769 = s_1770 - s_1777;
  assign s_1770 = s_1771;
  assign s_1771 = s_1772 | s_1776;
  assign s_1772 = s_1773 << s_1775;
  dq #(57, 1) dq_s_1773 (clk, s_1773, s_1774);
  assign s_1774 = s_1755?s_1758:s_1756;
  assign s_1775 = 1'd1;
  assign s_1776 = 1'd0;
  dq #(56, 6) dq_s_1777 (clk, s_1777, s_958);
  assign s_1778 = 1'd1;
  assign s_1779 = s_185 | s_1780;
  assign s_1780 = 1'd1;
  assign s_1781 = s_1782[56];
  assign s_1782 = s_1783 - s_1790;
  assign s_1783 = s_1784;
  assign s_1784 = s_1785 | s_1789;
  assign s_1785 = s_1786 << s_1788;
  dq #(57, 1) dq_s_1786 (clk, s_1786, s_1787);
  assign s_1787 = s_1768?s_1771:s_1769;
  assign s_1788 = 1'd1;
  assign s_1789 = 1'd0;
  dq #(56, 7) dq_s_1790 (clk, s_1790, s_958);
  assign s_1791 = 1'd1;
  assign s_1792 = s_182 | s_1793;
  assign s_1793 = 1'd1;
  assign s_1794 = s_1795[56];
  assign s_1795 = s_1796 - s_1803;
  assign s_1796 = s_1797;
  assign s_1797 = s_1798 | s_1802;
  assign s_1798 = s_1799 << s_1801;
  dq #(57, 1) dq_s_1799 (clk, s_1799, s_1800);
  assign s_1800 = s_1781?s_1784:s_1782;
  assign s_1801 = 1'd1;
  assign s_1802 = 1'd0;
  dq #(56, 8) dq_s_1803 (clk, s_1803, s_958);
  assign s_1804 = 1'd1;
  assign s_1805 = s_179 | s_1806;
  assign s_1806 = 1'd1;
  assign s_1807 = s_1808[56];
  assign s_1808 = s_1809 - s_1816;
  assign s_1809 = s_1810;
  assign s_1810 = s_1811 | s_1815;
  assign s_1811 = s_1812 << s_1814;
  dq #(57, 1) dq_s_1812 (clk, s_1812, s_1813);
  assign s_1813 = s_1794?s_1797:s_1795;
  assign s_1814 = 1'd1;
  assign s_1815 = 1'd0;
  dq #(56, 9) dq_s_1816 (clk, s_1816, s_958);
  assign s_1817 = 1'd1;
  assign s_1818 = s_176 | s_1819;
  assign s_1819 = 1'd1;
  assign s_1820 = s_1821[56];
  assign s_1821 = s_1822 - s_1829;
  assign s_1822 = s_1823;
  assign s_1823 = s_1824 | s_1828;
  assign s_1824 = s_1825 << s_1827;
  dq #(57, 1) dq_s_1825 (clk, s_1825, s_1826);
  assign s_1826 = s_1807?s_1810:s_1808;
  assign s_1827 = 1'd1;
  assign s_1828 = 1'd0;
  dq #(56, 10) dq_s_1829 (clk, s_1829, s_958);
  assign s_1830 = 1'd1;
  assign s_1831 = s_173 | s_1832;
  assign s_1832 = 1'd1;
  assign s_1833 = s_1834[56];
  assign s_1834 = s_1835 - s_1842;
  assign s_1835 = s_1836;
  assign s_1836 = s_1837 | s_1841;
  assign s_1837 = s_1838 << s_1840;
  dq #(57, 1) dq_s_1838 (clk, s_1838, s_1839);
  assign s_1839 = s_1820?s_1823:s_1821;
  assign s_1840 = 1'd1;
  assign s_1841 = 1'd0;
  dq #(56, 11) dq_s_1842 (clk, s_1842, s_958);
  assign s_1843 = 1'd1;
  assign s_1844 = s_170 | s_1845;
  assign s_1845 = 1'd1;
  assign s_1846 = s_1847[56];
  assign s_1847 = s_1848 - s_1855;
  assign s_1848 = s_1849;
  assign s_1849 = s_1850 | s_1854;
  assign s_1850 = s_1851 << s_1853;
  dq #(57, 1) dq_s_1851 (clk, s_1851, s_1852);
  assign s_1852 = s_1833?s_1836:s_1834;
  assign s_1853 = 1'd1;
  assign s_1854 = 1'd0;
  dq #(56, 12) dq_s_1855 (clk, s_1855, s_958);
  assign s_1856 = 1'd1;
  assign s_1857 = s_167 | s_1858;
  assign s_1858 = 1'd1;
  assign s_1859 = s_1860[56];
  assign s_1860 = s_1861 - s_1868;
  assign s_1861 = s_1862;
  assign s_1862 = s_1863 | s_1867;
  assign s_1863 = s_1864 << s_1866;
  dq #(57, 1) dq_s_1864 (clk, s_1864, s_1865);
  assign s_1865 = s_1846?s_1849:s_1847;
  assign s_1866 = 1'd1;
  assign s_1867 = 1'd0;
  dq #(56, 13) dq_s_1868 (clk, s_1868, s_958);
  assign s_1869 = 1'd1;
  assign s_1870 = s_164 | s_1871;
  assign s_1871 = 1'd1;
  assign s_1872 = s_1873[56];
  assign s_1873 = s_1874 - s_1881;
  assign s_1874 = s_1875;
  assign s_1875 = s_1876 | s_1880;
  assign s_1876 = s_1877 << s_1879;
  dq #(57, 1) dq_s_1877 (clk, s_1877, s_1878);
  assign s_1878 = s_1859?s_1862:s_1860;
  assign s_1879 = 1'd1;
  assign s_1880 = 1'd0;
  dq #(56, 14) dq_s_1881 (clk, s_1881, s_958);
  assign s_1882 = 1'd1;
  assign s_1883 = s_161 | s_1884;
  assign s_1884 = 1'd1;
  assign s_1885 = s_1886[56];
  assign s_1886 = s_1887 - s_1894;
  assign s_1887 = s_1888;
  assign s_1888 = s_1889 | s_1893;
  assign s_1889 = s_1890 << s_1892;
  dq #(57, 1) dq_s_1890 (clk, s_1890, s_1891);
  assign s_1891 = s_1872?s_1875:s_1873;
  assign s_1892 = 1'd1;
  assign s_1893 = 1'd0;
  dq #(56, 15) dq_s_1894 (clk, s_1894, s_958);
  assign s_1895 = 1'd1;
  assign s_1896 = s_158 | s_1897;
  assign s_1897 = 1'd1;
  assign s_1898 = s_1899[56];
  assign s_1899 = s_1900 - s_1907;
  assign s_1900 = s_1901;
  assign s_1901 = s_1902 | s_1906;
  assign s_1902 = s_1903 << s_1905;
  dq #(57, 1) dq_s_1903 (clk, s_1903, s_1904);
  assign s_1904 = s_1885?s_1888:s_1886;
  assign s_1905 = 1'd1;
  assign s_1906 = 1'd0;
  dq #(56, 16) dq_s_1907 (clk, s_1907, s_958);
  assign s_1908 = 1'd1;
  assign s_1909 = s_155 | s_1910;
  assign s_1910 = 1'd1;
  assign s_1911 = s_1912[56];
  assign s_1912 = s_1913 - s_1920;
  assign s_1913 = s_1914;
  assign s_1914 = s_1915 | s_1919;
  assign s_1915 = s_1916 << s_1918;
  dq #(57, 1) dq_s_1916 (clk, s_1916, s_1917);
  assign s_1917 = s_1898?s_1901:s_1899;
  assign s_1918 = 1'd1;
  assign s_1919 = 1'd0;
  dq #(56, 17) dq_s_1920 (clk, s_1920, s_958);
  assign s_1921 = 1'd1;
  assign s_1922 = s_152 | s_1923;
  assign s_1923 = 1'd1;
  assign s_1924 = s_1925[56];
  assign s_1925 = s_1926 - s_1933;
  assign s_1926 = s_1927;
  assign s_1927 = s_1928 | s_1932;
  assign s_1928 = s_1929 << s_1931;
  dq #(57, 1) dq_s_1929 (clk, s_1929, s_1930);
  assign s_1930 = s_1911?s_1914:s_1912;
  assign s_1931 = 1'd1;
  assign s_1932 = 1'd0;
  dq #(56, 18) dq_s_1933 (clk, s_1933, s_958);
  assign s_1934 = 1'd1;
  assign s_1935 = s_149 | s_1936;
  assign s_1936 = 1'd1;
  assign s_1937 = s_1938[56];
  assign s_1938 = s_1939 - s_1946;
  assign s_1939 = s_1940;
  assign s_1940 = s_1941 | s_1945;
  assign s_1941 = s_1942 << s_1944;
  dq #(57, 1) dq_s_1942 (clk, s_1942, s_1943);
  assign s_1943 = s_1924?s_1927:s_1925;
  assign s_1944 = 1'd1;
  assign s_1945 = 1'd0;
  dq #(56, 19) dq_s_1946 (clk, s_1946, s_958);
  assign s_1947 = 1'd1;
  assign s_1948 = s_146 | s_1949;
  assign s_1949 = 1'd1;
  assign s_1950 = s_1951[56];
  assign s_1951 = s_1952 - s_1959;
  assign s_1952 = s_1953;
  assign s_1953 = s_1954 | s_1958;
  assign s_1954 = s_1955 << s_1957;
  dq #(57, 1) dq_s_1955 (clk, s_1955, s_1956);
  assign s_1956 = s_1937?s_1940:s_1938;
  assign s_1957 = 1'd1;
  assign s_1958 = 1'd0;
  dq #(56, 20) dq_s_1959 (clk, s_1959, s_958);
  assign s_1960 = 1'd1;
  assign s_1961 = s_143 | s_1962;
  assign s_1962 = 1'd1;
  assign s_1963 = s_1964[56];
  assign s_1964 = s_1965 - s_1972;
  assign s_1965 = s_1966;
  assign s_1966 = s_1967 | s_1971;
  assign s_1967 = s_1968 << s_1970;
  dq #(57, 1) dq_s_1968 (clk, s_1968, s_1969);
  assign s_1969 = s_1950?s_1953:s_1951;
  assign s_1970 = 1'd1;
  assign s_1971 = 1'd0;
  dq #(56, 21) dq_s_1972 (clk, s_1972, s_958);
  assign s_1973 = 1'd1;
  assign s_1974 = s_140 | s_1975;
  assign s_1975 = 1'd1;
  assign s_1976 = s_1977[56];
  assign s_1977 = s_1978 - s_1985;
  assign s_1978 = s_1979;
  assign s_1979 = s_1980 | s_1984;
  assign s_1980 = s_1981 << s_1983;
  dq #(57, 1) dq_s_1981 (clk, s_1981, s_1982);
  assign s_1982 = s_1963?s_1966:s_1964;
  assign s_1983 = 1'd1;
  assign s_1984 = 1'd0;
  dq #(56, 22) dq_s_1985 (clk, s_1985, s_958);
  assign s_1986 = 1'd1;
  assign s_1987 = s_137 | s_1988;
  assign s_1988 = 1'd1;
  assign s_1989 = s_1990[56];
  assign s_1990 = s_1991 - s_1998;
  assign s_1991 = s_1992;
  assign s_1992 = s_1993 | s_1997;
  assign s_1993 = s_1994 << s_1996;
  dq #(57, 1) dq_s_1994 (clk, s_1994, s_1995);
  assign s_1995 = s_1976?s_1979:s_1977;
  assign s_1996 = 1'd1;
  assign s_1997 = 1'd0;
  dq #(56, 23) dq_s_1998 (clk, s_1998, s_958);
  assign s_1999 = 1'd1;
  assign s_2000 = s_134 | s_2001;
  assign s_2001 = 1'd1;
  assign s_2002 = s_2003[56];
  assign s_2003 = s_2004 - s_2011;
  assign s_2004 = s_2005;
  assign s_2005 = s_2006 | s_2010;
  assign s_2006 = s_2007 << s_2009;
  dq #(57, 1) dq_s_2007 (clk, s_2007, s_2008);
  assign s_2008 = s_1989?s_1992:s_1990;
  assign s_2009 = 1'd1;
  assign s_2010 = 1'd0;
  dq #(56, 24) dq_s_2011 (clk, s_2011, s_958);
  assign s_2012 = 1'd1;
  assign s_2013 = s_131 | s_2014;
  assign s_2014 = 1'd1;
  assign s_2015 = s_2016[56];
  assign s_2016 = s_2017 - s_2024;
  assign s_2017 = s_2018;
  assign s_2018 = s_2019 | s_2023;
  assign s_2019 = s_2020 << s_2022;
  dq #(57, 1) dq_s_2020 (clk, s_2020, s_2021);
  assign s_2021 = s_2002?s_2005:s_2003;
  assign s_2022 = 1'd1;
  assign s_2023 = 1'd0;
  dq #(56, 25) dq_s_2024 (clk, s_2024, s_958);
  assign s_2025 = 1'd1;
  assign s_2026 = s_128 | s_2027;
  assign s_2027 = 1'd1;
  assign s_2028 = s_2029[56];
  assign s_2029 = s_2030 - s_2037;
  assign s_2030 = s_2031;
  assign s_2031 = s_2032 | s_2036;
  assign s_2032 = s_2033 << s_2035;
  dq #(57, 1) dq_s_2033 (clk, s_2033, s_2034);
  assign s_2034 = s_2015?s_2018:s_2016;
  assign s_2035 = 1'd1;
  assign s_2036 = 1'd0;
  dq #(56, 26) dq_s_2037 (clk, s_2037, s_958);
  assign s_2038 = 1'd1;
  assign s_2039 = s_125 | s_2040;
  assign s_2040 = 1'd1;
  assign s_2041 = s_2042[56];
  assign s_2042 = s_2043 - s_2050;
  assign s_2043 = s_2044;
  assign s_2044 = s_2045 | s_2049;
  assign s_2045 = s_2046 << s_2048;
  dq #(57, 1) dq_s_2046 (clk, s_2046, s_2047);
  assign s_2047 = s_2028?s_2031:s_2029;
  assign s_2048 = 1'd1;
  assign s_2049 = 1'd0;
  dq #(56, 27) dq_s_2050 (clk, s_2050, s_958);
  assign s_2051 = 1'd1;
  assign s_2052 = s_122 | s_2053;
  assign s_2053 = 1'd1;
  assign s_2054 = s_2055[56];
  assign s_2055 = s_2056 - s_2063;
  assign s_2056 = s_2057;
  assign s_2057 = s_2058 | s_2062;
  assign s_2058 = s_2059 << s_2061;
  dq #(57, 1) dq_s_2059 (clk, s_2059, s_2060);
  assign s_2060 = s_2041?s_2044:s_2042;
  assign s_2061 = 1'd1;
  assign s_2062 = 1'd0;
  dq #(56, 28) dq_s_2063 (clk, s_2063, s_958);
  assign s_2064 = 1'd1;
  assign s_2065 = s_119 | s_2066;
  assign s_2066 = 1'd1;
  assign s_2067 = s_2068[56];
  assign s_2068 = s_2069 - s_2076;
  assign s_2069 = s_2070;
  assign s_2070 = s_2071 | s_2075;
  assign s_2071 = s_2072 << s_2074;
  dq #(57, 1) dq_s_2072 (clk, s_2072, s_2073);
  assign s_2073 = s_2054?s_2057:s_2055;
  assign s_2074 = 1'd1;
  assign s_2075 = 1'd0;
  dq #(56, 29) dq_s_2076 (clk, s_2076, s_958);
  assign s_2077 = 1'd1;
  assign s_2078 = s_116 | s_2079;
  assign s_2079 = 1'd1;
  assign s_2080 = s_2081[56];
  assign s_2081 = s_2082 - s_2089;
  assign s_2082 = s_2083;
  assign s_2083 = s_2084 | s_2088;
  assign s_2084 = s_2085 << s_2087;
  dq #(57, 1) dq_s_2085 (clk, s_2085, s_2086);
  assign s_2086 = s_2067?s_2070:s_2068;
  assign s_2087 = 1'd1;
  assign s_2088 = 1'd0;
  dq #(56, 30) dq_s_2089 (clk, s_2089, s_958);
  assign s_2090 = 1'd1;
  assign s_2091 = s_113 | s_2092;
  assign s_2092 = 1'd1;
  assign s_2093 = s_2094[56];
  assign s_2094 = s_2095 - s_2102;
  assign s_2095 = s_2096;
  assign s_2096 = s_2097 | s_2101;
  assign s_2097 = s_2098 << s_2100;
  dq #(57, 1) dq_s_2098 (clk, s_2098, s_2099);
  assign s_2099 = s_2080?s_2083:s_2081;
  assign s_2100 = 1'd1;
  assign s_2101 = 1'd0;
  dq #(56, 31) dq_s_2102 (clk, s_2102, s_958);
  assign s_2103 = 1'd1;
  assign s_2104 = s_110 | s_2105;
  assign s_2105 = 1'd1;
  assign s_2106 = s_2107[56];
  assign s_2107 = s_2108 - s_2115;
  assign s_2108 = s_2109;
  assign s_2109 = s_2110 | s_2114;
  assign s_2110 = s_2111 << s_2113;
  dq #(57, 1) dq_s_2111 (clk, s_2111, s_2112);
  assign s_2112 = s_2093?s_2096:s_2094;
  assign s_2113 = 1'd1;
  assign s_2114 = 1'd0;
  dq #(56, 32) dq_s_2115 (clk, s_2115, s_958);
  assign s_2116 = 1'd1;
  assign s_2117 = s_107 | s_2118;
  assign s_2118 = 1'd1;
  assign s_2119 = s_2120[56];
  assign s_2120 = s_2121 - s_2128;
  assign s_2121 = s_2122;
  assign s_2122 = s_2123 | s_2127;
  assign s_2123 = s_2124 << s_2126;
  dq #(57, 1) dq_s_2124 (clk, s_2124, s_2125);
  assign s_2125 = s_2106?s_2109:s_2107;
  assign s_2126 = 1'd1;
  assign s_2127 = 1'd0;
  dq #(56, 33) dq_s_2128 (clk, s_2128, s_958);
  assign s_2129 = 1'd1;
  assign s_2130 = s_104 | s_2131;
  assign s_2131 = 1'd1;
  assign s_2132 = s_2133[56];
  assign s_2133 = s_2134 - s_2141;
  assign s_2134 = s_2135;
  assign s_2135 = s_2136 | s_2140;
  assign s_2136 = s_2137 << s_2139;
  dq #(57, 1) dq_s_2137 (clk, s_2137, s_2138);
  assign s_2138 = s_2119?s_2122:s_2120;
  assign s_2139 = 1'd1;
  assign s_2140 = 1'd0;
  dq #(56, 34) dq_s_2141 (clk, s_2141, s_958);
  assign s_2142 = 1'd1;
  assign s_2143 = s_101 | s_2144;
  assign s_2144 = 1'd1;
  assign s_2145 = s_2146[56];
  assign s_2146 = s_2147 - s_2154;
  assign s_2147 = s_2148;
  assign s_2148 = s_2149 | s_2153;
  assign s_2149 = s_2150 << s_2152;
  dq #(57, 1) dq_s_2150 (clk, s_2150, s_2151);
  assign s_2151 = s_2132?s_2135:s_2133;
  assign s_2152 = 1'd1;
  assign s_2153 = 1'd0;
  dq #(56, 35) dq_s_2154 (clk, s_2154, s_958);
  assign s_2155 = 1'd1;
  assign s_2156 = s_98 | s_2157;
  assign s_2157 = 1'd1;
  assign s_2158 = s_2159[56];
  assign s_2159 = s_2160 - s_2167;
  assign s_2160 = s_2161;
  assign s_2161 = s_2162 | s_2166;
  assign s_2162 = s_2163 << s_2165;
  dq #(57, 1) dq_s_2163 (clk, s_2163, s_2164);
  assign s_2164 = s_2145?s_2148:s_2146;
  assign s_2165 = 1'd1;
  assign s_2166 = 1'd0;
  dq #(56, 36) dq_s_2167 (clk, s_2167, s_958);
  assign s_2168 = 1'd1;
  assign s_2169 = s_95 | s_2170;
  assign s_2170 = 1'd1;
  assign s_2171 = s_2172[56];
  assign s_2172 = s_2173 - s_2180;
  assign s_2173 = s_2174;
  assign s_2174 = s_2175 | s_2179;
  assign s_2175 = s_2176 << s_2178;
  dq #(57, 1) dq_s_2176 (clk, s_2176, s_2177);
  assign s_2177 = s_2158?s_2161:s_2159;
  assign s_2178 = 1'd1;
  assign s_2179 = 1'd0;
  dq #(56, 37) dq_s_2180 (clk, s_2180, s_958);
  assign s_2181 = 1'd1;
  assign s_2182 = s_92 | s_2183;
  assign s_2183 = 1'd1;
  assign s_2184 = s_2185[56];
  assign s_2185 = s_2186 - s_2193;
  assign s_2186 = s_2187;
  assign s_2187 = s_2188 | s_2192;
  assign s_2188 = s_2189 << s_2191;
  dq #(57, 1) dq_s_2189 (clk, s_2189, s_2190);
  assign s_2190 = s_2171?s_2174:s_2172;
  assign s_2191 = 1'd1;
  assign s_2192 = 1'd0;
  dq #(56, 38) dq_s_2193 (clk, s_2193, s_958);
  assign s_2194 = 1'd1;
  assign s_2195 = s_89 | s_2196;
  assign s_2196 = 1'd1;
  assign s_2197 = s_2198[56];
  assign s_2198 = s_2199 - s_2206;
  assign s_2199 = s_2200;
  assign s_2200 = s_2201 | s_2205;
  assign s_2201 = s_2202 << s_2204;
  dq #(57, 1) dq_s_2202 (clk, s_2202, s_2203);
  assign s_2203 = s_2184?s_2187:s_2185;
  assign s_2204 = 1'd1;
  assign s_2205 = 1'd0;
  dq #(56, 39) dq_s_2206 (clk, s_2206, s_958);
  assign s_2207 = 1'd1;
  assign s_2208 = s_86 | s_2209;
  assign s_2209 = 1'd1;
  assign s_2210 = s_2211[56];
  assign s_2211 = s_2212 - s_2219;
  assign s_2212 = s_2213;
  assign s_2213 = s_2214 | s_2218;
  assign s_2214 = s_2215 << s_2217;
  dq #(57, 1) dq_s_2215 (clk, s_2215, s_2216);
  assign s_2216 = s_2197?s_2200:s_2198;
  assign s_2217 = 1'd1;
  assign s_2218 = 1'd0;
  dq #(56, 40) dq_s_2219 (clk, s_2219, s_958);
  assign s_2220 = 1'd1;
  assign s_2221 = s_83 | s_2222;
  assign s_2222 = 1'd1;
  assign s_2223 = s_2224[56];
  assign s_2224 = s_2225 - s_2232;
  assign s_2225 = s_2226;
  assign s_2226 = s_2227 | s_2231;
  assign s_2227 = s_2228 << s_2230;
  dq #(57, 1) dq_s_2228 (clk, s_2228, s_2229);
  assign s_2229 = s_2210?s_2213:s_2211;
  assign s_2230 = 1'd1;
  assign s_2231 = 1'd0;
  dq #(56, 41) dq_s_2232 (clk, s_2232, s_958);
  assign s_2233 = 1'd1;
  assign s_2234 = s_80 | s_2235;
  assign s_2235 = 1'd1;
  assign s_2236 = s_2237[56];
  assign s_2237 = s_2238 - s_2245;
  assign s_2238 = s_2239;
  assign s_2239 = s_2240 | s_2244;
  assign s_2240 = s_2241 << s_2243;
  dq #(57, 1) dq_s_2241 (clk, s_2241, s_2242);
  assign s_2242 = s_2223?s_2226:s_2224;
  assign s_2243 = 1'd1;
  assign s_2244 = 1'd0;
  dq #(56, 42) dq_s_2245 (clk, s_2245, s_958);
  assign s_2246 = 1'd1;
  assign s_2247 = s_77 | s_2248;
  assign s_2248 = 1'd1;
  assign s_2249 = s_2250[56];
  assign s_2250 = s_2251 - s_2258;
  assign s_2251 = s_2252;
  assign s_2252 = s_2253 | s_2257;
  assign s_2253 = s_2254 << s_2256;
  dq #(57, 1) dq_s_2254 (clk, s_2254, s_2255);
  assign s_2255 = s_2236?s_2239:s_2237;
  assign s_2256 = 1'd1;
  assign s_2257 = 1'd0;
  dq #(56, 43) dq_s_2258 (clk, s_2258, s_958);
  assign s_2259 = 1'd1;
  assign s_2260 = s_74 | s_2261;
  assign s_2261 = 1'd1;
  assign s_2262 = s_2263[56];
  assign s_2263 = s_2264 - s_2271;
  assign s_2264 = s_2265;
  assign s_2265 = s_2266 | s_2270;
  assign s_2266 = s_2267 << s_2269;
  dq #(57, 1) dq_s_2267 (clk, s_2267, s_2268);
  assign s_2268 = s_2249?s_2252:s_2250;
  assign s_2269 = 1'd1;
  assign s_2270 = 1'd0;
  dq #(56, 44) dq_s_2271 (clk, s_2271, s_958);
  assign s_2272 = 1'd1;
  assign s_2273 = s_71 | s_2274;
  assign s_2274 = 1'd1;
  assign s_2275 = s_2276[56];
  assign s_2276 = s_2277 - s_2284;
  assign s_2277 = s_2278;
  assign s_2278 = s_2279 | s_2283;
  assign s_2279 = s_2280 << s_2282;
  dq #(57, 1) dq_s_2280 (clk, s_2280, s_2281);
  assign s_2281 = s_2262?s_2265:s_2263;
  assign s_2282 = 1'd1;
  assign s_2283 = 1'd0;
  dq #(56, 45) dq_s_2284 (clk, s_2284, s_958);
  assign s_2285 = 1'd1;
  assign s_2286 = s_68 | s_2287;
  assign s_2287 = 1'd1;
  assign s_2288 = s_2289[56];
  assign s_2289 = s_2290 - s_2297;
  assign s_2290 = s_2291;
  assign s_2291 = s_2292 | s_2296;
  assign s_2292 = s_2293 << s_2295;
  dq #(57, 1) dq_s_2293 (clk, s_2293, s_2294);
  assign s_2294 = s_2275?s_2278:s_2276;
  assign s_2295 = 1'd1;
  assign s_2296 = 1'd0;
  dq #(56, 46) dq_s_2297 (clk, s_2297, s_958);
  assign s_2298 = 1'd1;
  assign s_2299 = s_65 | s_2300;
  assign s_2300 = 1'd1;
  assign s_2301 = s_2302[56];
  assign s_2302 = s_2303 - s_2310;
  assign s_2303 = s_2304;
  assign s_2304 = s_2305 | s_2309;
  assign s_2305 = s_2306 << s_2308;
  dq #(57, 1) dq_s_2306 (clk, s_2306, s_2307);
  assign s_2307 = s_2288?s_2291:s_2289;
  assign s_2308 = 1'd1;
  assign s_2309 = 1'd0;
  dq #(56, 47) dq_s_2310 (clk, s_2310, s_958);
  assign s_2311 = 1'd1;
  assign s_2312 = s_62 | s_2313;
  assign s_2313 = 1'd1;
  assign s_2314 = s_2315[56];
  assign s_2315 = s_2316 - s_2323;
  assign s_2316 = s_2317;
  assign s_2317 = s_2318 | s_2322;
  assign s_2318 = s_2319 << s_2321;
  dq #(57, 1) dq_s_2319 (clk, s_2319, s_2320);
  assign s_2320 = s_2301?s_2304:s_2302;
  assign s_2321 = 1'd1;
  assign s_2322 = 1'd0;
  dq #(56, 48) dq_s_2323 (clk, s_2323, s_958);
  assign s_2324 = 1'd1;
  assign s_2325 = s_59 | s_2326;
  assign s_2326 = 1'd1;
  assign s_2327 = s_2328[56];
  assign s_2328 = s_2329 - s_2336;
  assign s_2329 = s_2330;
  assign s_2330 = s_2331 | s_2335;
  assign s_2331 = s_2332 << s_2334;
  dq #(57, 1) dq_s_2332 (clk, s_2332, s_2333);
  assign s_2333 = s_2314?s_2317:s_2315;
  assign s_2334 = 1'd1;
  assign s_2335 = 1'd0;
  dq #(56, 49) dq_s_2336 (clk, s_2336, s_958);
  assign s_2337 = 1'd1;
  assign s_2338 = s_56 | s_2339;
  assign s_2339 = 1'd1;
  assign s_2340 = s_2341[56];
  assign s_2341 = s_2342 - s_2349;
  assign s_2342 = s_2343;
  assign s_2343 = s_2344 | s_2348;
  assign s_2344 = s_2345 << s_2347;
  dq #(57, 1) dq_s_2345 (clk, s_2345, s_2346);
  assign s_2346 = s_2327?s_2330:s_2328;
  assign s_2347 = 1'd1;
  assign s_2348 = 1'd0;
  dq #(56, 50) dq_s_2349 (clk, s_2349, s_958);
  assign s_2350 = 1'd1;
  assign s_2351 = s_53 | s_2352;
  assign s_2352 = 1'd1;
  assign s_2353 = s_2354[56];
  assign s_2354 = s_2355 - s_2362;
  assign s_2355 = s_2356;
  assign s_2356 = s_2357 | s_2361;
  assign s_2357 = s_2358 << s_2360;
  dq #(57, 1) dq_s_2358 (clk, s_2358, s_2359);
  assign s_2359 = s_2340?s_2343:s_2341;
  assign s_2360 = 1'd1;
  assign s_2361 = 1'd0;
  dq #(56, 51) dq_s_2362 (clk, s_2362, s_958);
  assign s_2363 = 1'd1;
  assign s_2364 = s_50 | s_2365;
  assign s_2365 = 1'd1;
  assign s_2366 = s_2367[56];
  assign s_2367 = s_2368 - s_2375;
  assign s_2368 = s_2369;
  assign s_2369 = s_2370 | s_2374;
  assign s_2370 = s_2371 << s_2373;
  dq #(57, 1) dq_s_2371 (clk, s_2371, s_2372);
  assign s_2372 = s_2353?s_2356:s_2354;
  assign s_2373 = 1'd1;
  assign s_2374 = 1'd0;
  dq #(56, 52) dq_s_2375 (clk, s_2375, s_958);
  assign s_2376 = 1'd1;
  assign s_2377 = s_47 | s_2378;
  assign s_2378 = 1'd1;
  assign s_2379 = s_2380[56];
  assign s_2380 = s_2381 - s_2388;
  assign s_2381 = s_2382;
  assign s_2382 = s_2383 | s_2387;
  assign s_2383 = s_2384 << s_2386;
  dq #(57, 1) dq_s_2384 (clk, s_2384, s_2385);
  assign s_2385 = s_2366?s_2369:s_2367;
  assign s_2386 = 1'd1;
  assign s_2387 = 1'd0;
  dq #(56, 53) dq_s_2388 (clk, s_2388, s_958);
  assign s_2389 = 1'd1;
  assign s_2390 = s_44 | s_2391;
  assign s_2391 = 1'd1;
  assign s_2392 = s_2393[56];
  assign s_2393 = s_2394 - s_2401;
  assign s_2394 = s_2395;
  assign s_2395 = s_2396 | s_2400;
  assign s_2396 = s_2397 << s_2399;
  dq #(57, 1) dq_s_2397 (clk, s_2397, s_2398);
  assign s_2398 = s_2379?s_2382:s_2380;
  assign s_2399 = 1'd1;
  assign s_2400 = 1'd0;
  dq #(56, 54) dq_s_2401 (clk, s_2401, s_958);
  assign s_2402 = 1'd1;
  assign s_2403 = s_41 | s_2404;
  assign s_2404 = 1'd1;
  assign s_2405 = s_2406[56];
  assign s_2406 = s_2407 - s_2414;
  assign s_2407 = s_2408;
  assign s_2408 = s_2409 | s_2413;
  assign s_2409 = s_2410 << s_2412;
  dq #(57, 1) dq_s_2410 (clk, s_2410, s_2411);
  assign s_2411 = s_2392?s_2395:s_2393;
  assign s_2412 = 1'd1;
  assign s_2413 = 1'd0;
  dq #(56, 55) dq_s_2414 (clk, s_2414, s_958);
  dq #(13, 53) dq_s_2415 (clk, s_2415, s_2416);
  dq #(13, 1) dq_s_2416 (clk, s_2416, s_2417);
  assign s_2417 = s_2430?s_2418:s_2419;
  assign s_2418 = 1'd0;
  dq #(13, 1) dq_s_2419 (clk, s_2419, s_2420);
  assign s_2420 = s_2421 - s_2422;
  assign s_2421 = -13'd1022;
  dq #(13, 1) dq_s_2422 (clk, s_2422, s_2423);
  assign s_2423 = s_2424 - s_2427;
  dq #(13, 1) dq_s_2424 (clk, s_2424, s_2425);
  assign s_2425 = s_2426 - s_231;
  dq #(13, 2) dq_s_2426 (clk, s_2426, s_950);
  dq #(13, 1) dq_s_2427 (clk, s_2427, s_2428);
  assign s_2428 = s_2429 - s_973;
  dq #(13, 2) dq_s_2429 (clk, s_2429, s_1692);
  assign s_2430 = s_2419[12];
  dq #(13, 1) dq_s_2431 (clk, s_2431, s_2432);
  assign s_2432 = s_3148?s_2433:s_3142;
  dq #(7, 1) dq_s_2433 (clk, s_2433, s_2434);
  assign s_2434 = {s_2435,s_3136};
  assign s_2435 = s_2436 & s_2794;
  assign s_2436 = s_2437[5];
  assign s_2437 = {s_2438,s_2788};
  assign s_2438 = s_2439 & s_2622;
  assign s_2439 = s_2440[4];
  assign s_2440 = {s_2441,s_2616};
  assign s_2441 = s_2442 & s_2538;
  assign s_2442 = s_2443[3];
  assign s_2443 = {s_2444,s_2532};
  assign s_2444 = s_2445 & s_2498;
  assign s_2445 = s_2446[2];
  assign s_2446 = {s_2447,s_2492};
  assign s_2447 = s_2448 & s_2480;
  assign s_2448 = s_2449[1];
  assign s_2449 = {s_2450,s_2476};
  assign s_2450 = s_2451 & s_2474;
  assign s_2451 = ~s_2452;
  assign s_2452 = s_2453[1];
  assign s_2453 = s_2454[3:2];
  assign s_2454 = s_2455[7:4];
  assign s_2455 = s_2456[15:8];
  assign s_2456 = s_2457[31:16];
  assign s_2457 = s_2458[63:32];
  assign s_2458 = {s_2459,s_2473};
  assign s_2459 = {s_2460,s_2472};
  assign s_2460 = {s_2461,s_2471};
  assign s_2461 = {s_2462,s_2470};
  assign s_2462 = {s_2463,s_2469};
  assign s_2463 = {s_2464,s_2468};
  assign s_2464 = {s_2465,s_2467};
  assign s_2465 = {s_37,s_2466};
  assign s_2466 = 1'd1;
  assign s_2467 = 1'd1;
  assign s_2468 = 1'd1;
  assign s_2469 = 1'd1;
  assign s_2470 = 1'd1;
  assign s_2471 = 1'd1;
  assign s_2472 = 1'd1;
  assign s_2473 = 1'd1;
  assign s_2474 = ~s_2475;
  assign s_2475 = s_2453[0];
  assign s_2476 = s_2477 & s_2479;
  assign s_2477 = ~s_2478;
  assign s_2478 = s_2453[1];
  assign s_2479 = s_2453[0];
  assign s_2480 = s_2481[1];
  assign s_2481 = {s_2482,s_2488};
  assign s_2482 = s_2483 & s_2486;
  assign s_2483 = ~s_2484;
  assign s_2484 = s_2485[1];
  assign s_2485 = s_2454[1:0];
  assign s_2486 = ~s_2487;
  assign s_2487 = s_2485[0];
  assign s_2488 = s_2489 & s_2491;
  assign s_2489 = ~s_2490;
  assign s_2490 = s_2485[1];
  assign s_2491 = s_2485[0];
  assign s_2492 = {s_2493,s_2495};
  assign s_2493 = s_2448 & s_2494;
  assign s_2494 = ~s_2480;
  assign s_2495 = s_2448?s_2496:s_2497;
  assign s_2496 = s_2481[0:0];
  assign s_2497 = s_2449[0:0];
  assign s_2498 = s_2499[2];
  assign s_2499 = {s_2500,s_2526};
  assign s_2500 = s_2501 & s_2514;
  assign s_2501 = s_2502[1];
  assign s_2502 = {s_2503,s_2510};
  assign s_2503 = s_2504 & s_2508;
  assign s_2504 = ~s_2505;
  assign s_2505 = s_2506[1];
  assign s_2506 = s_2507[3:2];
  assign s_2507 = s_2455[3:0];
  assign s_2508 = ~s_2509;
  assign s_2509 = s_2506[0];
  assign s_2510 = s_2511 & s_2513;
  assign s_2511 = ~s_2512;
  assign s_2512 = s_2506[1];
  assign s_2513 = s_2506[0];
  assign s_2514 = s_2515[1];
  assign s_2515 = {s_2516,s_2522};
  assign s_2516 = s_2517 & s_2520;
  assign s_2517 = ~s_2518;
  assign s_2518 = s_2519[1];
  assign s_2519 = s_2507[1:0];
  assign s_2520 = ~s_2521;
  assign s_2521 = s_2519[0];
  assign s_2522 = s_2523 & s_2525;
  assign s_2523 = ~s_2524;
  assign s_2524 = s_2519[1];
  assign s_2525 = s_2519[0];
  assign s_2526 = {s_2527,s_2529};
  assign s_2527 = s_2501 & s_2528;
  assign s_2528 = ~s_2514;
  assign s_2529 = s_2501?s_2530:s_2531;
  assign s_2530 = s_2515[0:0];
  assign s_2531 = s_2502[0:0];
  assign s_2532 = {s_2533,s_2535};
  assign s_2533 = s_2445 & s_2534;
  assign s_2534 = ~s_2498;
  assign s_2535 = s_2445?s_2536:s_2537;
  assign s_2536 = s_2499[1:0];
  assign s_2537 = s_2446[1:0];
  assign s_2538 = s_2539[3];
  assign s_2539 = {s_2540,s_2610};
  assign s_2540 = s_2541 & s_2576;
  assign s_2541 = s_2542[2];
  assign s_2542 = {s_2543,s_2570};
  assign s_2543 = s_2544 & s_2558;
  assign s_2544 = s_2545[1];
  assign s_2545 = {s_2546,s_2554};
  assign s_2546 = s_2547 & s_2552;
  assign s_2547 = ~s_2548;
  assign s_2548 = s_2549[1];
  assign s_2549 = s_2550[3:2];
  assign s_2550 = s_2551[7:4];
  assign s_2551 = s_2456[7:0];
  assign s_2552 = ~s_2553;
  assign s_2553 = s_2549[0];
  assign s_2554 = s_2555 & s_2557;
  assign s_2555 = ~s_2556;
  assign s_2556 = s_2549[1];
  assign s_2557 = s_2549[0];
  assign s_2558 = s_2559[1];
  assign s_2559 = {s_2560,s_2566};
  assign s_2560 = s_2561 & s_2564;
  assign s_2561 = ~s_2562;
  assign s_2562 = s_2563[1];
  assign s_2563 = s_2550[1:0];
  assign s_2564 = ~s_2565;
  assign s_2565 = s_2563[0];
  assign s_2566 = s_2567 & s_2569;
  assign s_2567 = ~s_2568;
  assign s_2568 = s_2563[1];
  assign s_2569 = s_2563[0];
  assign s_2570 = {s_2571,s_2573};
  assign s_2571 = s_2544 & s_2572;
  assign s_2572 = ~s_2558;
  assign s_2573 = s_2544?s_2574:s_2575;
  assign s_2574 = s_2559[0:0];
  assign s_2575 = s_2545[0:0];
  assign s_2576 = s_2577[2];
  assign s_2577 = {s_2578,s_2604};
  assign s_2578 = s_2579 & s_2592;
  assign s_2579 = s_2580[1];
  assign s_2580 = {s_2581,s_2588};
  assign s_2581 = s_2582 & s_2586;
  assign s_2582 = ~s_2583;
  assign s_2583 = s_2584[1];
  assign s_2584 = s_2585[3:2];
  assign s_2585 = s_2551[3:0];
  assign s_2586 = ~s_2587;
  assign s_2587 = s_2584[0];
  assign s_2588 = s_2589 & s_2591;
  assign s_2589 = ~s_2590;
  assign s_2590 = s_2584[1];
  assign s_2591 = s_2584[0];
  assign s_2592 = s_2593[1];
  assign s_2593 = {s_2594,s_2600};
  assign s_2594 = s_2595 & s_2598;
  assign s_2595 = ~s_2596;
  assign s_2596 = s_2597[1];
  assign s_2597 = s_2585[1:0];
  assign s_2598 = ~s_2599;
  assign s_2599 = s_2597[0];
  assign s_2600 = s_2601 & s_2603;
  assign s_2601 = ~s_2602;
  assign s_2602 = s_2597[1];
  assign s_2603 = s_2597[0];
  assign s_2604 = {s_2605,s_2607};
  assign s_2605 = s_2579 & s_2606;
  assign s_2606 = ~s_2592;
  assign s_2607 = s_2579?s_2608:s_2609;
  assign s_2608 = s_2593[0:0];
  assign s_2609 = s_2580[0:0];
  assign s_2610 = {s_2611,s_2613};
  assign s_2611 = s_2541 & s_2612;
  assign s_2612 = ~s_2576;
  assign s_2613 = s_2541?s_2614:s_2615;
  assign s_2614 = s_2577[1:0];
  assign s_2615 = s_2542[1:0];
  assign s_2616 = {s_2617,s_2619};
  assign s_2617 = s_2442 & s_2618;
  assign s_2618 = ~s_2538;
  assign s_2619 = s_2442?s_2620:s_2621;
  assign s_2620 = s_2539[2:0];
  assign s_2621 = s_2443[2:0];
  assign s_2622 = s_2623[4];
  assign s_2623 = {s_2624,s_2782};
  assign s_2624 = s_2625 & s_2704;
  assign s_2625 = s_2626[3];
  assign s_2626 = {s_2627,s_2698};
  assign s_2627 = s_2628 & s_2664;
  assign s_2628 = s_2629[2];
  assign s_2629 = {s_2630,s_2658};
  assign s_2630 = s_2631 & s_2646;
  assign s_2631 = s_2632[1];
  assign s_2632 = {s_2633,s_2642};
  assign s_2633 = s_2634 & s_2640;
  assign s_2634 = ~s_2635;
  assign s_2635 = s_2636[1];
  assign s_2636 = s_2637[3:2];
  assign s_2637 = s_2638[7:4];
  assign s_2638 = s_2639[15:8];
  assign s_2639 = s_2457[15:0];
  assign s_2640 = ~s_2641;
  assign s_2641 = s_2636[0];
  assign s_2642 = s_2643 & s_2645;
  assign s_2643 = ~s_2644;
  assign s_2644 = s_2636[1];
  assign s_2645 = s_2636[0];
  assign s_2646 = s_2647[1];
  assign s_2647 = {s_2648,s_2654};
  assign s_2648 = s_2649 & s_2652;
  assign s_2649 = ~s_2650;
  assign s_2650 = s_2651[1];
  assign s_2651 = s_2637[1:0];
  assign s_2652 = ~s_2653;
  assign s_2653 = s_2651[0];
  assign s_2654 = s_2655 & s_2657;
  assign s_2655 = ~s_2656;
  assign s_2656 = s_2651[1];
  assign s_2657 = s_2651[0];
  assign s_2658 = {s_2659,s_2661};
  assign s_2659 = s_2631 & s_2660;
  assign s_2660 = ~s_2646;
  assign s_2661 = s_2631?s_2662:s_2663;
  assign s_2662 = s_2647[0:0];
  assign s_2663 = s_2632[0:0];
  assign s_2664 = s_2665[2];
  assign s_2665 = {s_2666,s_2692};
  assign s_2666 = s_2667 & s_2680;
  assign s_2667 = s_2668[1];
  assign s_2668 = {s_2669,s_2676};
  assign s_2669 = s_2670 & s_2674;
  assign s_2670 = ~s_2671;
  assign s_2671 = s_2672[1];
  assign s_2672 = s_2673[3:2];
  assign s_2673 = s_2638[3:0];
  assign s_2674 = ~s_2675;
  assign s_2675 = s_2672[0];
  assign s_2676 = s_2677 & s_2679;
  assign s_2677 = ~s_2678;
  assign s_2678 = s_2672[1];
  assign s_2679 = s_2672[0];
  assign s_2680 = s_2681[1];
  assign s_2681 = {s_2682,s_2688};
  assign s_2682 = s_2683 & s_2686;
  assign s_2683 = ~s_2684;
  assign s_2684 = s_2685[1];
  assign s_2685 = s_2673[1:0];
  assign s_2686 = ~s_2687;
  assign s_2687 = s_2685[0];
  assign s_2688 = s_2689 & s_2691;
  assign s_2689 = ~s_2690;
  assign s_2690 = s_2685[1];
  assign s_2691 = s_2685[0];
  assign s_2692 = {s_2693,s_2695};
  assign s_2693 = s_2667 & s_2694;
  assign s_2694 = ~s_2680;
  assign s_2695 = s_2667?s_2696:s_2697;
  assign s_2696 = s_2681[0:0];
  assign s_2697 = s_2668[0:0];
  assign s_2698 = {s_2699,s_2701};
  assign s_2699 = s_2628 & s_2700;
  assign s_2700 = ~s_2664;
  assign s_2701 = s_2628?s_2702:s_2703;
  assign s_2702 = s_2665[1:0];
  assign s_2703 = s_2629[1:0];
  assign s_2704 = s_2705[3];
  assign s_2705 = {s_2706,s_2776};
  assign s_2706 = s_2707 & s_2742;
  assign s_2707 = s_2708[2];
  assign s_2708 = {s_2709,s_2736};
  assign s_2709 = s_2710 & s_2724;
  assign s_2710 = s_2711[1];
  assign s_2711 = {s_2712,s_2720};
  assign s_2712 = s_2713 & s_2718;
  assign s_2713 = ~s_2714;
  assign s_2714 = s_2715[1];
  assign s_2715 = s_2716[3:2];
  assign s_2716 = s_2717[7:4];
  assign s_2717 = s_2639[7:0];
  assign s_2718 = ~s_2719;
  assign s_2719 = s_2715[0];
  assign s_2720 = s_2721 & s_2723;
  assign s_2721 = ~s_2722;
  assign s_2722 = s_2715[1];
  assign s_2723 = s_2715[0];
  assign s_2724 = s_2725[1];
  assign s_2725 = {s_2726,s_2732};
  assign s_2726 = s_2727 & s_2730;
  assign s_2727 = ~s_2728;
  assign s_2728 = s_2729[1];
  assign s_2729 = s_2716[1:0];
  assign s_2730 = ~s_2731;
  assign s_2731 = s_2729[0];
  assign s_2732 = s_2733 & s_2735;
  assign s_2733 = ~s_2734;
  assign s_2734 = s_2729[1];
  assign s_2735 = s_2729[0];
  assign s_2736 = {s_2737,s_2739};
  assign s_2737 = s_2710 & s_2738;
  assign s_2738 = ~s_2724;
  assign s_2739 = s_2710?s_2740:s_2741;
  assign s_2740 = s_2725[0:0];
  assign s_2741 = s_2711[0:0];
  assign s_2742 = s_2743[2];
  assign s_2743 = {s_2744,s_2770};
  assign s_2744 = s_2745 & s_2758;
  assign s_2745 = s_2746[1];
  assign s_2746 = {s_2747,s_2754};
  assign s_2747 = s_2748 & s_2752;
  assign s_2748 = ~s_2749;
  assign s_2749 = s_2750[1];
  assign s_2750 = s_2751[3:2];
  assign s_2751 = s_2717[3:0];
  assign s_2752 = ~s_2753;
  assign s_2753 = s_2750[0];
  assign s_2754 = s_2755 & s_2757;
  assign s_2755 = ~s_2756;
  assign s_2756 = s_2750[1];
  assign s_2757 = s_2750[0];
  assign s_2758 = s_2759[1];
  assign s_2759 = {s_2760,s_2766};
  assign s_2760 = s_2761 & s_2764;
  assign s_2761 = ~s_2762;
  assign s_2762 = s_2763[1];
  assign s_2763 = s_2751[1:0];
  assign s_2764 = ~s_2765;
  assign s_2765 = s_2763[0];
  assign s_2766 = s_2767 & s_2769;
  assign s_2767 = ~s_2768;
  assign s_2768 = s_2763[1];
  assign s_2769 = s_2763[0];
  assign s_2770 = {s_2771,s_2773};
  assign s_2771 = s_2745 & s_2772;
  assign s_2772 = ~s_2758;
  assign s_2773 = s_2745?s_2774:s_2775;
  assign s_2774 = s_2759[0:0];
  assign s_2775 = s_2746[0:0];
  assign s_2776 = {s_2777,s_2779};
  assign s_2777 = s_2707 & s_2778;
  assign s_2778 = ~s_2742;
  assign s_2779 = s_2707?s_2780:s_2781;
  assign s_2780 = s_2743[1:0];
  assign s_2781 = s_2708[1:0];
  assign s_2782 = {s_2783,s_2785};
  assign s_2783 = s_2625 & s_2784;
  assign s_2784 = ~s_2704;
  assign s_2785 = s_2625?s_2786:s_2787;
  assign s_2786 = s_2705[2:0];
  assign s_2787 = s_2626[2:0];
  assign s_2788 = {s_2789,s_2791};
  assign s_2789 = s_2439 & s_2790;
  assign s_2790 = ~s_2622;
  assign s_2791 = s_2439?s_2792:s_2793;
  assign s_2792 = s_2623[3:0];
  assign s_2793 = s_2440[3:0];
  assign s_2794 = s_2795[5];
  assign s_2795 = {s_2796,s_3130};
  assign s_2796 = s_2797 & s_2964;
  assign s_2797 = s_2798[4];
  assign s_2798 = {s_2799,s_2958};
  assign s_2799 = s_2800 & s_2880;
  assign s_2800 = s_2801[3];
  assign s_2801 = {s_2802,s_2874};
  assign s_2802 = s_2803 & s_2840;
  assign s_2803 = s_2804[2];
  assign s_2804 = {s_2805,s_2834};
  assign s_2805 = s_2806 & s_2822;
  assign s_2806 = s_2807[1];
  assign s_2807 = {s_2808,s_2818};
  assign s_2808 = s_2809 & s_2816;
  assign s_2809 = ~s_2810;
  assign s_2810 = s_2811[1];
  assign s_2811 = s_2812[3:2];
  assign s_2812 = s_2813[7:4];
  assign s_2813 = s_2814[15:8];
  assign s_2814 = s_2815[31:16];
  assign s_2815 = s_2458[31:0];
  assign s_2816 = ~s_2817;
  assign s_2817 = s_2811[0];
  assign s_2818 = s_2819 & s_2821;
  assign s_2819 = ~s_2820;
  assign s_2820 = s_2811[1];
  assign s_2821 = s_2811[0];
  assign s_2822 = s_2823[1];
  assign s_2823 = {s_2824,s_2830};
  assign s_2824 = s_2825 & s_2828;
  assign s_2825 = ~s_2826;
  assign s_2826 = s_2827[1];
  assign s_2827 = s_2812[1:0];
  assign s_2828 = ~s_2829;
  assign s_2829 = s_2827[0];
  assign s_2830 = s_2831 & s_2833;
  assign s_2831 = ~s_2832;
  assign s_2832 = s_2827[1];
  assign s_2833 = s_2827[0];
  assign s_2834 = {s_2835,s_2837};
  assign s_2835 = s_2806 & s_2836;
  assign s_2836 = ~s_2822;
  assign s_2837 = s_2806?s_2838:s_2839;
  assign s_2838 = s_2823[0:0];
  assign s_2839 = s_2807[0:0];
  assign s_2840 = s_2841[2];
  assign s_2841 = {s_2842,s_2868};
  assign s_2842 = s_2843 & s_2856;
  assign s_2843 = s_2844[1];
  assign s_2844 = {s_2845,s_2852};
  assign s_2845 = s_2846 & s_2850;
  assign s_2846 = ~s_2847;
  assign s_2847 = s_2848[1];
  assign s_2848 = s_2849[3:2];
  assign s_2849 = s_2813[3:0];
  assign s_2850 = ~s_2851;
  assign s_2851 = s_2848[0];
  assign s_2852 = s_2853 & s_2855;
  assign s_2853 = ~s_2854;
  assign s_2854 = s_2848[1];
  assign s_2855 = s_2848[0];
  assign s_2856 = s_2857[1];
  assign s_2857 = {s_2858,s_2864};
  assign s_2858 = s_2859 & s_2862;
  assign s_2859 = ~s_2860;
  assign s_2860 = s_2861[1];
  assign s_2861 = s_2849[1:0];
  assign s_2862 = ~s_2863;
  assign s_2863 = s_2861[0];
  assign s_2864 = s_2865 & s_2867;
  assign s_2865 = ~s_2866;
  assign s_2866 = s_2861[1];
  assign s_2867 = s_2861[0];
  assign s_2868 = {s_2869,s_2871};
  assign s_2869 = s_2843 & s_2870;
  assign s_2870 = ~s_2856;
  assign s_2871 = s_2843?s_2872:s_2873;
  assign s_2872 = s_2857[0:0];
  assign s_2873 = s_2844[0:0];
  assign s_2874 = {s_2875,s_2877};
  assign s_2875 = s_2803 & s_2876;
  assign s_2876 = ~s_2840;
  assign s_2877 = s_2803?s_2878:s_2879;
  assign s_2878 = s_2841[1:0];
  assign s_2879 = s_2804[1:0];
  assign s_2880 = s_2881[3];
  assign s_2881 = {s_2882,s_2952};
  assign s_2882 = s_2883 & s_2918;
  assign s_2883 = s_2884[2];
  assign s_2884 = {s_2885,s_2912};
  assign s_2885 = s_2886 & s_2900;
  assign s_2886 = s_2887[1];
  assign s_2887 = {s_2888,s_2896};
  assign s_2888 = s_2889 & s_2894;
  assign s_2889 = ~s_2890;
  assign s_2890 = s_2891[1];
  assign s_2891 = s_2892[3:2];
  assign s_2892 = s_2893[7:4];
  assign s_2893 = s_2814[7:0];
  assign s_2894 = ~s_2895;
  assign s_2895 = s_2891[0];
  assign s_2896 = s_2897 & s_2899;
  assign s_2897 = ~s_2898;
  assign s_2898 = s_2891[1];
  assign s_2899 = s_2891[0];
  assign s_2900 = s_2901[1];
  assign s_2901 = {s_2902,s_2908};
  assign s_2902 = s_2903 & s_2906;
  assign s_2903 = ~s_2904;
  assign s_2904 = s_2905[1];
  assign s_2905 = s_2892[1:0];
  assign s_2906 = ~s_2907;
  assign s_2907 = s_2905[0];
  assign s_2908 = s_2909 & s_2911;
  assign s_2909 = ~s_2910;
  assign s_2910 = s_2905[1];
  assign s_2911 = s_2905[0];
  assign s_2912 = {s_2913,s_2915};
  assign s_2913 = s_2886 & s_2914;
  assign s_2914 = ~s_2900;
  assign s_2915 = s_2886?s_2916:s_2917;
  assign s_2916 = s_2901[0:0];
  assign s_2917 = s_2887[0:0];
  assign s_2918 = s_2919[2];
  assign s_2919 = {s_2920,s_2946};
  assign s_2920 = s_2921 & s_2934;
  assign s_2921 = s_2922[1];
  assign s_2922 = {s_2923,s_2930};
  assign s_2923 = s_2924 & s_2928;
  assign s_2924 = ~s_2925;
  assign s_2925 = s_2926[1];
  assign s_2926 = s_2927[3:2];
  assign s_2927 = s_2893[3:0];
  assign s_2928 = ~s_2929;
  assign s_2929 = s_2926[0];
  assign s_2930 = s_2931 & s_2933;
  assign s_2931 = ~s_2932;
  assign s_2932 = s_2926[1];
  assign s_2933 = s_2926[0];
  assign s_2934 = s_2935[1];
  assign s_2935 = {s_2936,s_2942};
  assign s_2936 = s_2937 & s_2940;
  assign s_2937 = ~s_2938;
  assign s_2938 = s_2939[1];
  assign s_2939 = s_2927[1:0];
  assign s_2940 = ~s_2941;
  assign s_2941 = s_2939[0];
  assign s_2942 = s_2943 & s_2945;
  assign s_2943 = ~s_2944;
  assign s_2944 = s_2939[1];
  assign s_2945 = s_2939[0];
  assign s_2946 = {s_2947,s_2949};
  assign s_2947 = s_2921 & s_2948;
  assign s_2948 = ~s_2934;
  assign s_2949 = s_2921?s_2950:s_2951;
  assign s_2950 = s_2935[0:0];
  assign s_2951 = s_2922[0:0];
  assign s_2952 = {s_2953,s_2955};
  assign s_2953 = s_2883 & s_2954;
  assign s_2954 = ~s_2918;
  assign s_2955 = s_2883?s_2956:s_2957;
  assign s_2956 = s_2919[1:0];
  assign s_2957 = s_2884[1:0];
  assign s_2958 = {s_2959,s_2961};
  assign s_2959 = s_2800 & s_2960;
  assign s_2960 = ~s_2880;
  assign s_2961 = s_2800?s_2962:s_2963;
  assign s_2962 = s_2881[2:0];
  assign s_2963 = s_2801[2:0];
  assign s_2964 = s_2965[4];
  assign s_2965 = {s_2966,s_3124};
  assign s_2966 = s_2967 & s_3046;
  assign s_2967 = s_2968[3];
  assign s_2968 = {s_2969,s_3040};
  assign s_2969 = s_2970 & s_3006;
  assign s_2970 = s_2971[2];
  assign s_2971 = {s_2972,s_3000};
  assign s_2972 = s_2973 & s_2988;
  assign s_2973 = s_2974[1];
  assign s_2974 = {s_2975,s_2984};
  assign s_2975 = s_2976 & s_2982;
  assign s_2976 = ~s_2977;
  assign s_2977 = s_2978[1];
  assign s_2978 = s_2979[3:2];
  assign s_2979 = s_2980[7:4];
  assign s_2980 = s_2981[15:8];
  assign s_2981 = s_2815[15:0];
  assign s_2982 = ~s_2983;
  assign s_2983 = s_2978[0];
  assign s_2984 = s_2985 & s_2987;
  assign s_2985 = ~s_2986;
  assign s_2986 = s_2978[1];
  assign s_2987 = s_2978[0];
  assign s_2988 = s_2989[1];
  assign s_2989 = {s_2990,s_2996};
  assign s_2990 = s_2991 & s_2994;
  assign s_2991 = ~s_2992;
  assign s_2992 = s_2993[1];
  assign s_2993 = s_2979[1:0];
  assign s_2994 = ~s_2995;
  assign s_2995 = s_2993[0];
  assign s_2996 = s_2997 & s_2999;
  assign s_2997 = ~s_2998;
  assign s_2998 = s_2993[1];
  assign s_2999 = s_2993[0];
  assign s_3000 = {s_3001,s_3003};
  assign s_3001 = s_2973 & s_3002;
  assign s_3002 = ~s_2988;
  assign s_3003 = s_2973?s_3004:s_3005;
  assign s_3004 = s_2989[0:0];
  assign s_3005 = s_2974[0:0];
  assign s_3006 = s_3007[2];
  assign s_3007 = {s_3008,s_3034};
  assign s_3008 = s_3009 & s_3022;
  assign s_3009 = s_3010[1];
  assign s_3010 = {s_3011,s_3018};
  assign s_3011 = s_3012 & s_3016;
  assign s_3012 = ~s_3013;
  assign s_3013 = s_3014[1];
  assign s_3014 = s_3015[3:2];
  assign s_3015 = s_2980[3:0];
  assign s_3016 = ~s_3017;
  assign s_3017 = s_3014[0];
  assign s_3018 = s_3019 & s_3021;
  assign s_3019 = ~s_3020;
  assign s_3020 = s_3014[1];
  assign s_3021 = s_3014[0];
  assign s_3022 = s_3023[1];
  assign s_3023 = {s_3024,s_3030};
  assign s_3024 = s_3025 & s_3028;
  assign s_3025 = ~s_3026;
  assign s_3026 = s_3027[1];
  assign s_3027 = s_3015[1:0];
  assign s_3028 = ~s_3029;
  assign s_3029 = s_3027[0];
  assign s_3030 = s_3031 & s_3033;
  assign s_3031 = ~s_3032;
  assign s_3032 = s_3027[1];
  assign s_3033 = s_3027[0];
  assign s_3034 = {s_3035,s_3037};
  assign s_3035 = s_3009 & s_3036;
  assign s_3036 = ~s_3022;
  assign s_3037 = s_3009?s_3038:s_3039;
  assign s_3038 = s_3023[0:0];
  assign s_3039 = s_3010[0:0];
  assign s_3040 = {s_3041,s_3043};
  assign s_3041 = s_2970 & s_3042;
  assign s_3042 = ~s_3006;
  assign s_3043 = s_2970?s_3044:s_3045;
  assign s_3044 = s_3007[1:0];
  assign s_3045 = s_2971[1:0];
  assign s_3046 = s_3047[3];
  assign s_3047 = {s_3048,s_3118};
  assign s_3048 = s_3049 & s_3084;
  assign s_3049 = s_3050[2];
  assign s_3050 = {s_3051,s_3078};
  assign s_3051 = s_3052 & s_3066;
  assign s_3052 = s_3053[1];
  assign s_3053 = {s_3054,s_3062};
  assign s_3054 = s_3055 & s_3060;
  assign s_3055 = ~s_3056;
  assign s_3056 = s_3057[1];
  assign s_3057 = s_3058[3:2];
  assign s_3058 = s_3059[7:4];
  assign s_3059 = s_2981[7:0];
  assign s_3060 = ~s_3061;
  assign s_3061 = s_3057[0];
  assign s_3062 = s_3063 & s_3065;
  assign s_3063 = ~s_3064;
  assign s_3064 = s_3057[1];
  assign s_3065 = s_3057[0];
  assign s_3066 = s_3067[1];
  assign s_3067 = {s_3068,s_3074};
  assign s_3068 = s_3069 & s_3072;
  assign s_3069 = ~s_3070;
  assign s_3070 = s_3071[1];
  assign s_3071 = s_3058[1:0];
  assign s_3072 = ~s_3073;
  assign s_3073 = s_3071[0];
  assign s_3074 = s_3075 & s_3077;
  assign s_3075 = ~s_3076;
  assign s_3076 = s_3071[1];
  assign s_3077 = s_3071[0];
  assign s_3078 = {s_3079,s_3081};
  assign s_3079 = s_3052 & s_3080;
  assign s_3080 = ~s_3066;
  assign s_3081 = s_3052?s_3082:s_3083;
  assign s_3082 = s_3067[0:0];
  assign s_3083 = s_3053[0:0];
  assign s_3084 = s_3085[2];
  assign s_3085 = {s_3086,s_3112};
  assign s_3086 = s_3087 & s_3100;
  assign s_3087 = s_3088[1];
  assign s_3088 = {s_3089,s_3096};
  assign s_3089 = s_3090 & s_3094;
  assign s_3090 = ~s_3091;
  assign s_3091 = s_3092[1];
  assign s_3092 = s_3093[3:2];
  assign s_3093 = s_3059[3:0];
  assign s_3094 = ~s_3095;
  assign s_3095 = s_3092[0];
  assign s_3096 = s_3097 & s_3099;
  assign s_3097 = ~s_3098;
  assign s_3098 = s_3092[1];
  assign s_3099 = s_3092[0];
  assign s_3100 = s_3101[1];
  assign s_3101 = {s_3102,s_3108};
  assign s_3102 = s_3103 & s_3106;
  assign s_3103 = ~s_3104;
  assign s_3104 = s_3105[1];
  assign s_3105 = s_3093[1:0];
  assign s_3106 = ~s_3107;
  assign s_3107 = s_3105[0];
  assign s_3108 = s_3109 & s_3111;
  assign s_3109 = ~s_3110;
  assign s_3110 = s_3105[1];
  assign s_3111 = s_3105[0];
  assign s_3112 = {s_3113,s_3115};
  assign s_3113 = s_3087 & s_3114;
  assign s_3114 = ~s_3100;
  assign s_3115 = s_3087?s_3116:s_3117;
  assign s_3116 = s_3101[0:0];
  assign s_3117 = s_3088[0:0];
  assign s_3118 = {s_3119,s_3121};
  assign s_3119 = s_3049 & s_3120;
  assign s_3120 = ~s_3084;
  assign s_3121 = s_3049?s_3122:s_3123;
  assign s_3122 = s_3085[1:0];
  assign s_3123 = s_3050[1:0];
  assign s_3124 = {s_3125,s_3127};
  assign s_3125 = s_2967 & s_3126;
  assign s_3126 = ~s_3046;
  assign s_3127 = s_2967?s_3128:s_3129;
  assign s_3128 = s_3047[2:0];
  assign s_3129 = s_2968[2:0];
  assign s_3130 = {s_3131,s_3133};
  assign s_3131 = s_2797 & s_3132;
  assign s_3132 = ~s_2964;
  assign s_3133 = s_2797?s_3134:s_3135;
  assign s_3134 = s_2965[3:0];
  assign s_3135 = s_2798[3:0];
  assign s_3136 = {s_3137,s_3139};
  assign s_3137 = s_2436 & s_3138;
  assign s_3138 = ~s_2794;
  assign s_3139 = s_2436?s_3140:s_3141;
  assign s_3140 = s_2795[4:0];
  assign s_3141 = s_2437[4:0];
  dq #(13, 54) dq_s_3142 (clk, s_3142, s_3143);
  assign s_3143 = s_3144 - s_3147;
  dq #(13, 1) dq_s_3144 (clk, s_3144, s_3145);
  assign s_3145 = s_3146 + s_2416;
  dq #(13, 2) dq_s_3146 (clk, s_3146, s_2422);
  assign s_3147 = -13'd1022;
  assign s_3148 = s_3149 <= s_3150;
  assign s_3149 = s_2433;
  dq #(13, 54) dq_s_3150 (clk, s_3150, s_3143);
  assign s_3151 = 2'd3;
  assign s_3152 = 1'd1;
  dq #(53, 1) dq_s_3153 (clk, s_3153, s_32);
  assign s_3154 = s_3155 & s_3157;
  dq #(1, 1) dq_s_3155 (clk, s_3155, s_3156);
  assign s_3156 = s_34[2];
  assign s_3157 = s_3158 | s_3169;
  assign s_3158 = s_3159 | s_3161;
  dq #(1, 1) dq_s_3159 (clk, s_3159, s_3160);
  assign s_3160 = s_34[1];
  dq #(1, 1) dq_s_3161 (clk, s_3161, s_3162);
  assign s_3162 = s_3163 | s_3164;
  assign s_3163 = s_34[0];
  dq #(1, 4) dq_s_3164 (clk, s_3164, s_3165);
  assign s_3165 = s_3166 != s_3168;
  dq #(57, 1) dq_s_3166 (clk, s_3166, s_3167);
  assign s_3167 = s_2405?s_2408:s_2406;
  assign s_3168 = 1'd0;
  dq #(1, 1) dq_s_3169 (clk, s_3169, s_3170);
  assign s_3170 = s_32[0];
  assign s_3171 = s_28[52:0];
  assign s_3172 = s_28[53];
  dq #(1, 65) dq_s_3173 (clk, s_3173, s_3174);
  assign s_3174 = s_3175 & s_3177;
  assign s_3175 = s_968 == s_3176;
  assign s_3176 = 11'd1024;
  assign s_3177 = s_972 == s_3178;
  assign s_3178 = 52'd0;
  assign s_3179 = {s_3180,s_3191};
  assign s_3180 = {s_3181,s_3182};
  dq #(1, 65) dq_s_3181 (clk, s_3181, s_3);
  assign s_3182 = s_3183 + s_3190;
  assign s_3183 = s_3184[10:0];
  dq #(13, 1) dq_s_3184 (clk, s_3184, s_3185);
  assign s_3185 = s_3186 + s_3172;
  dq #(13, 1) dq_s_3186 (clk, s_3186, s_3187);
  dq #(13, 1) dq_s_3187 (clk, s_3187, s_3188);
  assign s_3188 = s_3189 - s_2431;
  dq #(13, 55) dq_s_3189 (clk, s_3189, s_3144);
  assign s_3190 = 10'd1023;
  assign s_3191 = s_23[51:0];
  assign s_3192 = s_3193 & s_3195;
  assign s_3193 = s_3183 == s_3194;
  assign s_3194 = -11'd1022;
  assign s_3195 = ~s_3196;
  assign s_3196 = s_23[52];
  assign s_3197 = s_23 == s_3198;
  assign s_3198 = 53'd0;
  assign s_3199 = s_3215?s_3200:s_3201;
  assign s_3200 = 1'd0;
  assign s_3201 = s_3202 | s_3211;
  assign s_3202 = s_3203 | s_3205;
  assign s_3203 = $signed(s_3184) > $signed(s_3204);
  assign s_3204 = 12'd1023;
  dq #(1, 65) dq_s_3205 (clk, s_3205, s_3206);
  assign s_3206 = s_3207 & s_3209;
  assign s_3207 = s_226 == s_3208;
  assign s_3208 = 11'd1024;
  assign s_3209 = s_230 == s_3210;
  assign s_3210 = 52'd0;
  dq #(1, 61) dq_s_3211 (clk, s_3211, s_3212);
  dq #(1, 1) dq_s_3212 (clk, s_3212, s_3213);
  assign s_3213 = s_958 == s_3214;
  assign s_3214 = 1'd0;
  dq #(1, 65) dq_s_3215 (clk, s_3215, s_3174);
  dq #(1, 65) dq_s_3216 (clk, s_3216, s_3217);
  assign s_3217 = s_3218 | s_3229;
  assign s_3218 = s_3219 | s_3224;
  assign s_3219 = s_3220 & s_3222;
  assign s_3220 = s_226 == s_3221;
  assign s_3221 = 11'd1024;
  assign s_3222 = s_230 != s_3223;
  assign s_3223 = 52'd0;
  assign s_3224 = s_3225 & s_3227;
  assign s_3225 = s_968 == s_3226;
  assign s_3226 = 11'd1024;
  assign s_3227 = s_972 != s_3228;
  assign s_3228 = 52'd0;
  assign s_3229 = s_3206 & s_3174;
  assign double_div_z = s_0;
endmodule
