module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module mul(clk, mul_a, mul_b, mul_z);
  input clk;
  input [31:0] mul_a;
  input [31:0] mul_b;
  output [31:0] mul_z;
  wire [31:0] s_0;
  wire [31:0] s_1;
  wire [31:0] s_2;
  wire [0:0] s_3;
  wire [0:0] s_4;
  wire [31:0] s_5;
  wire [0:0] s_6;
  wire [31:0] s_7;
  wire [30:0] s_8;
  wire [31:0] s_9;
  wire [31:0] s_10;
  wire [31:0] s_11;
  wire [30:0] s_12;
  wire [31:0] s_13;
  wire [31:0] s_14;
  wire [31:0] s_15;
  wire [30:0] s_16;
  wire [31:0] s_17;
  wire [31:0] s_18;
  wire [8:0] s_19;
  wire [8:0] s_20;
  wire [7:0] s_21;
  wire [22:0] s_22;
  wire [23:0] s_23;
  wire [23:0] s_24;
  wire [23:0] s_25;
  wire [24:0] s_26;
  wire [24:0] s_27;
  wire [24:0] s_28;
  wire [24:0] s_29;
  wire [23:0] s_30;
  wire [47:0] s_31;
  wire [47:0] s_32;
  wire [47:0] s_33;
  wire [47:0] s_34;
  wire [47:0] s_35;
  wire [47:0] s_36;
  wire [50:0] s_37;
  wire [16:0] s_38;
  wire [33:0] s_39;
  wire [33:0] s_40;
  wire [33:0] s_41;
  wire [33:0] s_42;
  wire [33:0] s_43;
  wire [16:0] s_44;
  wire [33:0] s_45;
  wire [23:0] s_46;
  wire [0:0] s_47;
  wire [0:0] s_48;
  wire [0:0] s_49;
  wire [0:0] s_50;
  wire [7:0] s_51;
  wire [7:0] s_52;
  wire [6:0] s_53;
  wire [7:0] s_54;
  wire [22:0] s_55;
  wire [16:0] s_56;
  wire [33:0] s_57;
  wire [23:0] s_58;
  wire [0:0] s_59;
  wire [0:0] s_60;
  wire [0:0] s_61;
  wire [0:0] s_62;
  wire [7:0] s_63;
  wire [7:0] s_64;
  wire [6:0] s_65;
  wire [7:0] s_66;
  wire [22:0] s_67;
  wire [33:0] s_68;
  wire [33:0] s_69;
  wire [33:0] s_70;
  wire [33:0] s_71;
  wire [33:0] s_72;
  wire [33:0] s_73;
  wire [16:0] s_74;
  wire [33:0] s_75;
  wire [33:0] s_76;
  wire [33:0] s_77;
  wire [33:0] s_78;
  wire [16:0] s_79;
  wire [33:0] s_80;
  wire [33:0] s_81;
  wire [33:0] s_82;
  wire [4:0] s_83;
  wire [4:0] s_84;
  wire [33:0] s_85;
  wire [33:0] s_86;
  wire [16:0] s_87;
  wire [16:0] s_88;
  wire [16:0] s_89;
  wire [9:0] s_90;
  wire [9:0] s_91;
  wire [0:0] s_92;
  wire [9:0] s_93;
  wire [9:0] s_94;
  wire [9:0] s_95;
  wire [9:0] s_96;
  wire [9:0] s_97;
  wire [7:0] s_98;
  wire [7:0] s_99;
  wire [9:0] s_100;
  wire [7:0] s_101;
  wire [7:0] s_102;
  wire [0:0] s_103;
  wire [0:0] s_104;
  wire [9:0] s_105;
  wire [9:0] s_106;
  wire [6:0] s_107;
  wire [6:0] s_108;
  wire [0:0] s_109;
  wire [0:0] s_110;
  wire [5:0] s_111;
  wire [0:0] s_112;
  wire [0:0] s_113;
  wire [4:0] s_114;
  wire [0:0] s_115;
  wire [0:0] s_116;
  wire [3:0] s_117;
  wire [0:0] s_118;
  wire [0:0] s_119;
  wire [2:0] s_120;
  wire [0:0] s_121;
  wire [0:0] s_122;
  wire [1:0] s_123;
  wire [0:0] s_124;
  wire [0:0] s_125;
  wire [0:0] s_126;
  wire [1:0] s_127;
  wire [3:0] s_128;
  wire [7:0] s_129;
  wire [15:0] s_130;
  wire [31:0] s_131;
  wire [63:0] s_132;
  wire [62:0] s_133;
  wire [61:0] s_134;
  wire [60:0] s_135;
  wire [59:0] s_136;
  wire [58:0] s_137;
  wire [57:0] s_138;
  wire [56:0] s_139;
  wire [55:0] s_140;
  wire [54:0] s_141;
  wire [53:0] s_142;
  wire [52:0] s_143;
  wire [51:0] s_144;
  wire [50:0] s_145;
  wire [49:0] s_146;
  wire [48:0] s_147;
  wire [0:0] s_148;
  wire [0:0] s_149;
  wire [0:0] s_150;
  wire [0:0] s_151;
  wire [0:0] s_152;
  wire [0:0] s_153;
  wire [0:0] s_154;
  wire [0:0] s_155;
  wire [0:0] s_156;
  wire [0:0] s_157;
  wire [0:0] s_158;
  wire [0:0] s_159;
  wire [0:0] s_160;
  wire [0:0] s_161;
  wire [0:0] s_162;
  wire [0:0] s_163;
  wire [0:0] s_164;
  wire [0:0] s_165;
  wire [0:0] s_166;
  wire [0:0] s_167;
  wire [0:0] s_168;
  wire [0:0] s_169;
  wire [0:0] s_170;
  wire [1:0] s_171;
  wire [0:0] s_172;
  wire [0:0] s_173;
  wire [0:0] s_174;
  wire [1:0] s_175;
  wire [0:0] s_176;
  wire [0:0] s_177;
  wire [0:0] s_178;
  wire [0:0] s_179;
  wire [0:0] s_180;
  wire [0:0] s_181;
  wire [1:0] s_182;
  wire [0:0] s_183;
  wire [0:0] s_184;
  wire [0:0] s_185;
  wire [0:0] s_186;
  wire [0:0] s_187;
  wire [0:0] s_188;
  wire [2:0] s_189;
  wire [0:0] s_190;
  wire [0:0] s_191;
  wire [1:0] s_192;
  wire [0:0] s_193;
  wire [0:0] s_194;
  wire [0:0] s_195;
  wire [1:0] s_196;
  wire [3:0] s_197;
  wire [0:0] s_198;
  wire [0:0] s_199;
  wire [0:0] s_200;
  wire [0:0] s_201;
  wire [0:0] s_202;
  wire [0:0] s_203;
  wire [0:0] s_204;
  wire [1:0] s_205;
  wire [0:0] s_206;
  wire [0:0] s_207;
  wire [0:0] s_208;
  wire [1:0] s_209;
  wire [0:0] s_210;
  wire [0:0] s_211;
  wire [0:0] s_212;
  wire [0:0] s_213;
  wire [0:0] s_214;
  wire [0:0] s_215;
  wire [1:0] s_216;
  wire [0:0] s_217;
  wire [0:0] s_218;
  wire [0:0] s_219;
  wire [0:0] s_220;
  wire [0:0] s_221;
  wire [2:0] s_222;
  wire [0:0] s_223;
  wire [0:0] s_224;
  wire [1:0] s_225;
  wire [1:0] s_226;
  wire [1:0] s_227;
  wire [0:0] s_228;
  wire [3:0] s_229;
  wire [0:0] s_230;
  wire [0:0] s_231;
  wire [2:0] s_232;
  wire [0:0] s_233;
  wire [0:0] s_234;
  wire [1:0] s_235;
  wire [0:0] s_236;
  wire [0:0] s_237;
  wire [0:0] s_238;
  wire [1:0] s_239;
  wire [3:0] s_240;
  wire [7:0] s_241;
  wire [0:0] s_242;
  wire [0:0] s_243;
  wire [0:0] s_244;
  wire [0:0] s_245;
  wire [0:0] s_246;
  wire [0:0] s_247;
  wire [0:0] s_248;
  wire [1:0] s_249;
  wire [0:0] s_250;
  wire [0:0] s_251;
  wire [0:0] s_252;
  wire [1:0] s_253;
  wire [0:0] s_254;
  wire [0:0] s_255;
  wire [0:0] s_256;
  wire [0:0] s_257;
  wire [0:0] s_258;
  wire [0:0] s_259;
  wire [1:0] s_260;
  wire [0:0] s_261;
  wire [0:0] s_262;
  wire [0:0] s_263;
  wire [0:0] s_264;
  wire [0:0] s_265;
  wire [0:0] s_266;
  wire [2:0] s_267;
  wire [0:0] s_268;
  wire [0:0] s_269;
  wire [1:0] s_270;
  wire [0:0] s_271;
  wire [0:0] s_272;
  wire [0:0] s_273;
  wire [1:0] s_274;
  wire [3:0] s_275;
  wire [0:0] s_276;
  wire [0:0] s_277;
  wire [0:0] s_278;
  wire [0:0] s_279;
  wire [0:0] s_280;
  wire [0:0] s_281;
  wire [0:0] s_282;
  wire [1:0] s_283;
  wire [0:0] s_284;
  wire [0:0] s_285;
  wire [0:0] s_286;
  wire [1:0] s_287;
  wire [0:0] s_288;
  wire [0:0] s_289;
  wire [0:0] s_290;
  wire [0:0] s_291;
  wire [0:0] s_292;
  wire [0:0] s_293;
  wire [1:0] s_294;
  wire [0:0] s_295;
  wire [0:0] s_296;
  wire [0:0] s_297;
  wire [0:0] s_298;
  wire [0:0] s_299;
  wire [2:0] s_300;
  wire [0:0] s_301;
  wire [0:0] s_302;
  wire [1:0] s_303;
  wire [1:0] s_304;
  wire [1:0] s_305;
  wire [3:0] s_306;
  wire [0:0] s_307;
  wire [0:0] s_308;
  wire [2:0] s_309;
  wire [2:0] s_310;
  wire [2:0] s_311;
  wire [0:0] s_312;
  wire [4:0] s_313;
  wire [0:0] s_314;
  wire [0:0] s_315;
  wire [3:0] s_316;
  wire [0:0] s_317;
  wire [0:0] s_318;
  wire [2:0] s_319;
  wire [0:0] s_320;
  wire [0:0] s_321;
  wire [1:0] s_322;
  wire [0:0] s_323;
  wire [0:0] s_324;
  wire [0:0] s_325;
  wire [1:0] s_326;
  wire [3:0] s_327;
  wire [7:0] s_328;
  wire [15:0] s_329;
  wire [0:0] s_330;
  wire [0:0] s_331;
  wire [0:0] s_332;
  wire [0:0] s_333;
  wire [0:0] s_334;
  wire [0:0] s_335;
  wire [0:0] s_336;
  wire [1:0] s_337;
  wire [0:0] s_338;
  wire [0:0] s_339;
  wire [0:0] s_340;
  wire [1:0] s_341;
  wire [0:0] s_342;
  wire [0:0] s_343;
  wire [0:0] s_344;
  wire [0:0] s_345;
  wire [0:0] s_346;
  wire [0:0] s_347;
  wire [1:0] s_348;
  wire [0:0] s_349;
  wire [0:0] s_350;
  wire [0:0] s_351;
  wire [0:0] s_352;
  wire [0:0] s_353;
  wire [0:0] s_354;
  wire [2:0] s_355;
  wire [0:0] s_356;
  wire [0:0] s_357;
  wire [1:0] s_358;
  wire [0:0] s_359;
  wire [0:0] s_360;
  wire [0:0] s_361;
  wire [1:0] s_362;
  wire [3:0] s_363;
  wire [0:0] s_364;
  wire [0:0] s_365;
  wire [0:0] s_366;
  wire [0:0] s_367;
  wire [0:0] s_368;
  wire [0:0] s_369;
  wire [0:0] s_370;
  wire [1:0] s_371;
  wire [0:0] s_372;
  wire [0:0] s_373;
  wire [0:0] s_374;
  wire [1:0] s_375;
  wire [0:0] s_376;
  wire [0:0] s_377;
  wire [0:0] s_378;
  wire [0:0] s_379;
  wire [0:0] s_380;
  wire [0:0] s_381;
  wire [1:0] s_382;
  wire [0:0] s_383;
  wire [0:0] s_384;
  wire [0:0] s_385;
  wire [0:0] s_386;
  wire [0:0] s_387;
  wire [2:0] s_388;
  wire [0:0] s_389;
  wire [0:0] s_390;
  wire [1:0] s_391;
  wire [1:0] s_392;
  wire [1:0] s_393;
  wire [0:0] s_394;
  wire [3:0] s_395;
  wire [0:0] s_396;
  wire [0:0] s_397;
  wire [2:0] s_398;
  wire [0:0] s_399;
  wire [0:0] s_400;
  wire [1:0] s_401;
  wire [0:0] s_402;
  wire [0:0] s_403;
  wire [0:0] s_404;
  wire [1:0] s_405;
  wire [3:0] s_406;
  wire [7:0] s_407;
  wire [0:0] s_408;
  wire [0:0] s_409;
  wire [0:0] s_410;
  wire [0:0] s_411;
  wire [0:0] s_412;
  wire [0:0] s_413;
  wire [0:0] s_414;
  wire [1:0] s_415;
  wire [0:0] s_416;
  wire [0:0] s_417;
  wire [0:0] s_418;
  wire [1:0] s_419;
  wire [0:0] s_420;
  wire [0:0] s_421;
  wire [0:0] s_422;
  wire [0:0] s_423;
  wire [0:0] s_424;
  wire [0:0] s_425;
  wire [1:0] s_426;
  wire [0:0] s_427;
  wire [0:0] s_428;
  wire [0:0] s_429;
  wire [0:0] s_430;
  wire [0:0] s_431;
  wire [0:0] s_432;
  wire [2:0] s_433;
  wire [0:0] s_434;
  wire [0:0] s_435;
  wire [1:0] s_436;
  wire [0:0] s_437;
  wire [0:0] s_438;
  wire [0:0] s_439;
  wire [1:0] s_440;
  wire [3:0] s_441;
  wire [0:0] s_442;
  wire [0:0] s_443;
  wire [0:0] s_444;
  wire [0:0] s_445;
  wire [0:0] s_446;
  wire [0:0] s_447;
  wire [0:0] s_448;
  wire [1:0] s_449;
  wire [0:0] s_450;
  wire [0:0] s_451;
  wire [0:0] s_452;
  wire [1:0] s_453;
  wire [0:0] s_454;
  wire [0:0] s_455;
  wire [0:0] s_456;
  wire [0:0] s_457;
  wire [0:0] s_458;
  wire [0:0] s_459;
  wire [1:0] s_460;
  wire [0:0] s_461;
  wire [0:0] s_462;
  wire [0:0] s_463;
  wire [0:0] s_464;
  wire [0:0] s_465;
  wire [2:0] s_466;
  wire [0:0] s_467;
  wire [0:0] s_468;
  wire [1:0] s_469;
  wire [1:0] s_470;
  wire [1:0] s_471;
  wire [3:0] s_472;
  wire [0:0] s_473;
  wire [0:0] s_474;
  wire [2:0] s_475;
  wire [2:0] s_476;
  wire [2:0] s_477;
  wire [4:0] s_478;
  wire [0:0] s_479;
  wire [0:0] s_480;
  wire [3:0] s_481;
  wire [3:0] s_482;
  wire [3:0] s_483;
  wire [0:0] s_484;
  wire [5:0] s_485;
  wire [0:0] s_486;
  wire [0:0] s_487;
  wire [4:0] s_488;
  wire [0:0] s_489;
  wire [0:0] s_490;
  wire [3:0] s_491;
  wire [0:0] s_492;
  wire [0:0] s_493;
  wire [2:0] s_494;
  wire [0:0] s_495;
  wire [0:0] s_496;
  wire [1:0] s_497;
  wire [0:0] s_498;
  wire [0:0] s_499;
  wire [0:0] s_500;
  wire [1:0] s_501;
  wire [3:0] s_502;
  wire [7:0] s_503;
  wire [15:0] s_504;
  wire [31:0] s_505;
  wire [0:0] s_506;
  wire [0:0] s_507;
  wire [0:0] s_508;
  wire [0:0] s_509;
  wire [0:0] s_510;
  wire [0:0] s_511;
  wire [0:0] s_512;
  wire [1:0] s_513;
  wire [0:0] s_514;
  wire [0:0] s_515;
  wire [0:0] s_516;
  wire [1:0] s_517;
  wire [0:0] s_518;
  wire [0:0] s_519;
  wire [0:0] s_520;
  wire [0:0] s_521;
  wire [0:0] s_522;
  wire [0:0] s_523;
  wire [1:0] s_524;
  wire [0:0] s_525;
  wire [0:0] s_526;
  wire [0:0] s_527;
  wire [0:0] s_528;
  wire [0:0] s_529;
  wire [0:0] s_530;
  wire [2:0] s_531;
  wire [0:0] s_532;
  wire [0:0] s_533;
  wire [1:0] s_534;
  wire [0:0] s_535;
  wire [0:0] s_536;
  wire [0:0] s_537;
  wire [1:0] s_538;
  wire [3:0] s_539;
  wire [0:0] s_540;
  wire [0:0] s_541;
  wire [0:0] s_542;
  wire [0:0] s_543;
  wire [0:0] s_544;
  wire [0:0] s_545;
  wire [0:0] s_546;
  wire [1:0] s_547;
  wire [0:0] s_548;
  wire [0:0] s_549;
  wire [0:0] s_550;
  wire [1:0] s_551;
  wire [0:0] s_552;
  wire [0:0] s_553;
  wire [0:0] s_554;
  wire [0:0] s_555;
  wire [0:0] s_556;
  wire [0:0] s_557;
  wire [1:0] s_558;
  wire [0:0] s_559;
  wire [0:0] s_560;
  wire [0:0] s_561;
  wire [0:0] s_562;
  wire [0:0] s_563;
  wire [2:0] s_564;
  wire [0:0] s_565;
  wire [0:0] s_566;
  wire [1:0] s_567;
  wire [1:0] s_568;
  wire [1:0] s_569;
  wire [0:0] s_570;
  wire [3:0] s_571;
  wire [0:0] s_572;
  wire [0:0] s_573;
  wire [2:0] s_574;
  wire [0:0] s_575;
  wire [0:0] s_576;
  wire [1:0] s_577;
  wire [0:0] s_578;
  wire [0:0] s_579;
  wire [0:0] s_580;
  wire [1:0] s_581;
  wire [3:0] s_582;
  wire [7:0] s_583;
  wire [0:0] s_584;
  wire [0:0] s_585;
  wire [0:0] s_586;
  wire [0:0] s_587;
  wire [0:0] s_588;
  wire [0:0] s_589;
  wire [0:0] s_590;
  wire [1:0] s_591;
  wire [0:0] s_592;
  wire [0:0] s_593;
  wire [0:0] s_594;
  wire [1:0] s_595;
  wire [0:0] s_596;
  wire [0:0] s_597;
  wire [0:0] s_598;
  wire [0:0] s_599;
  wire [0:0] s_600;
  wire [0:0] s_601;
  wire [1:0] s_602;
  wire [0:0] s_603;
  wire [0:0] s_604;
  wire [0:0] s_605;
  wire [0:0] s_606;
  wire [0:0] s_607;
  wire [0:0] s_608;
  wire [2:0] s_609;
  wire [0:0] s_610;
  wire [0:0] s_611;
  wire [1:0] s_612;
  wire [0:0] s_613;
  wire [0:0] s_614;
  wire [0:0] s_615;
  wire [1:0] s_616;
  wire [3:0] s_617;
  wire [0:0] s_618;
  wire [0:0] s_619;
  wire [0:0] s_620;
  wire [0:0] s_621;
  wire [0:0] s_622;
  wire [0:0] s_623;
  wire [0:0] s_624;
  wire [1:0] s_625;
  wire [0:0] s_626;
  wire [0:0] s_627;
  wire [0:0] s_628;
  wire [1:0] s_629;
  wire [0:0] s_630;
  wire [0:0] s_631;
  wire [0:0] s_632;
  wire [0:0] s_633;
  wire [0:0] s_634;
  wire [0:0] s_635;
  wire [1:0] s_636;
  wire [0:0] s_637;
  wire [0:0] s_638;
  wire [0:0] s_639;
  wire [0:0] s_640;
  wire [0:0] s_641;
  wire [2:0] s_642;
  wire [0:0] s_643;
  wire [0:0] s_644;
  wire [1:0] s_645;
  wire [1:0] s_646;
  wire [1:0] s_647;
  wire [3:0] s_648;
  wire [0:0] s_649;
  wire [0:0] s_650;
  wire [2:0] s_651;
  wire [2:0] s_652;
  wire [2:0] s_653;
  wire [0:0] s_654;
  wire [4:0] s_655;
  wire [0:0] s_656;
  wire [0:0] s_657;
  wire [3:0] s_658;
  wire [0:0] s_659;
  wire [0:0] s_660;
  wire [2:0] s_661;
  wire [0:0] s_662;
  wire [0:0] s_663;
  wire [1:0] s_664;
  wire [0:0] s_665;
  wire [0:0] s_666;
  wire [0:0] s_667;
  wire [1:0] s_668;
  wire [3:0] s_669;
  wire [7:0] s_670;
  wire [15:0] s_671;
  wire [0:0] s_672;
  wire [0:0] s_673;
  wire [0:0] s_674;
  wire [0:0] s_675;
  wire [0:0] s_676;
  wire [0:0] s_677;
  wire [0:0] s_678;
  wire [1:0] s_679;
  wire [0:0] s_680;
  wire [0:0] s_681;
  wire [0:0] s_682;
  wire [1:0] s_683;
  wire [0:0] s_684;
  wire [0:0] s_685;
  wire [0:0] s_686;
  wire [0:0] s_687;
  wire [0:0] s_688;
  wire [0:0] s_689;
  wire [1:0] s_690;
  wire [0:0] s_691;
  wire [0:0] s_692;
  wire [0:0] s_693;
  wire [0:0] s_694;
  wire [0:0] s_695;
  wire [0:0] s_696;
  wire [2:0] s_697;
  wire [0:0] s_698;
  wire [0:0] s_699;
  wire [1:0] s_700;
  wire [0:0] s_701;
  wire [0:0] s_702;
  wire [0:0] s_703;
  wire [1:0] s_704;
  wire [3:0] s_705;
  wire [0:0] s_706;
  wire [0:0] s_707;
  wire [0:0] s_708;
  wire [0:0] s_709;
  wire [0:0] s_710;
  wire [0:0] s_711;
  wire [0:0] s_712;
  wire [1:0] s_713;
  wire [0:0] s_714;
  wire [0:0] s_715;
  wire [0:0] s_716;
  wire [1:0] s_717;
  wire [0:0] s_718;
  wire [0:0] s_719;
  wire [0:0] s_720;
  wire [0:0] s_721;
  wire [0:0] s_722;
  wire [0:0] s_723;
  wire [1:0] s_724;
  wire [0:0] s_725;
  wire [0:0] s_726;
  wire [0:0] s_727;
  wire [0:0] s_728;
  wire [0:0] s_729;
  wire [2:0] s_730;
  wire [0:0] s_731;
  wire [0:0] s_732;
  wire [1:0] s_733;
  wire [1:0] s_734;
  wire [1:0] s_735;
  wire [0:0] s_736;
  wire [3:0] s_737;
  wire [0:0] s_738;
  wire [0:0] s_739;
  wire [2:0] s_740;
  wire [0:0] s_741;
  wire [0:0] s_742;
  wire [1:0] s_743;
  wire [0:0] s_744;
  wire [0:0] s_745;
  wire [0:0] s_746;
  wire [1:0] s_747;
  wire [3:0] s_748;
  wire [7:0] s_749;
  wire [0:0] s_750;
  wire [0:0] s_751;
  wire [0:0] s_752;
  wire [0:0] s_753;
  wire [0:0] s_754;
  wire [0:0] s_755;
  wire [0:0] s_756;
  wire [1:0] s_757;
  wire [0:0] s_758;
  wire [0:0] s_759;
  wire [0:0] s_760;
  wire [1:0] s_761;
  wire [0:0] s_762;
  wire [0:0] s_763;
  wire [0:0] s_764;
  wire [0:0] s_765;
  wire [0:0] s_766;
  wire [0:0] s_767;
  wire [1:0] s_768;
  wire [0:0] s_769;
  wire [0:0] s_770;
  wire [0:0] s_771;
  wire [0:0] s_772;
  wire [0:0] s_773;
  wire [0:0] s_774;
  wire [2:0] s_775;
  wire [0:0] s_776;
  wire [0:0] s_777;
  wire [1:0] s_778;
  wire [0:0] s_779;
  wire [0:0] s_780;
  wire [0:0] s_781;
  wire [1:0] s_782;
  wire [3:0] s_783;
  wire [0:0] s_784;
  wire [0:0] s_785;
  wire [0:0] s_786;
  wire [0:0] s_787;
  wire [0:0] s_788;
  wire [0:0] s_789;
  wire [0:0] s_790;
  wire [1:0] s_791;
  wire [0:0] s_792;
  wire [0:0] s_793;
  wire [0:0] s_794;
  wire [1:0] s_795;
  wire [0:0] s_796;
  wire [0:0] s_797;
  wire [0:0] s_798;
  wire [0:0] s_799;
  wire [0:0] s_800;
  wire [0:0] s_801;
  wire [1:0] s_802;
  wire [0:0] s_803;
  wire [0:0] s_804;
  wire [0:0] s_805;
  wire [0:0] s_806;
  wire [0:0] s_807;
  wire [2:0] s_808;
  wire [0:0] s_809;
  wire [0:0] s_810;
  wire [1:0] s_811;
  wire [1:0] s_812;
  wire [1:0] s_813;
  wire [3:0] s_814;
  wire [0:0] s_815;
  wire [0:0] s_816;
  wire [2:0] s_817;
  wire [2:0] s_818;
  wire [2:0] s_819;
  wire [4:0] s_820;
  wire [0:0] s_821;
  wire [0:0] s_822;
  wire [3:0] s_823;
  wire [3:0] s_824;
  wire [3:0] s_825;
  wire [5:0] s_826;
  wire [0:0] s_827;
  wire [0:0] s_828;
  wire [4:0] s_829;
  wire [4:0] s_830;
  wire [4:0] s_831;
  wire [9:0] s_832;
  wire [9:0] s_833;
  wire [9:0] s_834;
  wire [9:0] s_835;
  wire [9:0] s_836;
  wire [0:0] s_837;
  wire [9:0] s_838;
  wire [9:0] s_839;
  wire [0:0] s_840;
  wire [23:0] s_841;
  wire [0:0] s_842;
  wire [0:0] s_843;
  wire [0:0] s_844;
  wire [0:0] s_845;
  wire [0:0] s_846;
  wire [0:0] s_847;
  wire [0:0] s_848;
  wire [0:0] s_849;
  wire [0:0] s_850;
  wire [21:0] s_851;
  wire [23:0] s_852;
  wire [0:0] s_853;
  wire [0:0] s_854;
  wire [23:0] s_855;
  wire [0:0] s_856;
  wire [31:0] s_857;
  wire [8:0] s_858;
  wire [0:0] s_859;
  wire [7:0] s_860;
  wire [7:0] s_861;
  wire [9:0] s_862;
  wire [9:0] s_863;
  wire [9:0] s_864;
  wire [9:0] s_865;
  wire [9:0] s_866;
  wire [9:0] s_867;
  wire [6:0] s_868;
  wire [22:0] s_869;
  wire [0:0] s_870;
  wire [0:0] s_871;
  wire [7:0] s_872;
  wire [0:0] s_873;
  wire [0:0] s_874;
  wire [0:0] s_875;
  wire [23:0] s_876;
  wire [0:0] s_877;
  wire [0:0] s_878;
  wire [0:0] s_879;
  wire [8:0] s_880;
  wire [0:0] s_881;
  wire [0:0] s_882;
  wire [0:0] s_883;
  wire [7:0] s_884;
  wire [0:0] s_885;
  wire [22:0] s_886;
  wire [0:0] s_887;
  wire [0:0] s_888;
  wire [0:0] s_889;
  wire [7:0] s_890;
  wire [0:0] s_891;
  wire [22:0] s_892;
  wire [0:0] s_893;
  wire [0:0] s_894;
  wire [0:0] s_895;
  wire [0:0] s_896;
  wire [7:0] s_897;
  wire [0:0] s_898;
  wire [22:0] s_899;
  wire [0:0] s_900;
  wire [0:0] s_901;
  wire [7:0] s_902;
  wire [0:0] s_903;
  wire [22:0] s_904;

  assign s_0 = s_893?s_1:s_9;
  dq #(32, 9) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_8};
  assign s_3 = s_4 ^ s_6;
  assign s_4 = s_5[31];
  assign s_5 = mul_a;
  assign s_6 = s_7[31];
  assign s_7 = mul_b;
  assign s_8 = 31'd2143289344;
  assign s_9 = s_877?s_10:s_13;
  dq #(32, 9) dq_s_10 (clk, s_10, s_11);
  assign s_11 = {s_3,s_12};
  assign s_12 = 31'd2139095040;
  assign s_13 = s_875?s_14:s_17;
  dq #(32, 9) dq_s_14 (clk, s_14, s_15);
  assign s_15 = {s_3,s_16};
  assign s_16 = 31'd0;
  assign s_17 = s_870?s_18:s_857;
  assign s_18 = {s_19,s_22};
  dq #(9, 9) dq_s_19 (clk, s_19, s_20);
  assign s_20 = {s_3,s_21};
  assign s_21 = 8'd0;
  assign s_22 = s_23[22:0];
  dq #(24, 1) dq_s_23 (clk, s_23, s_24);
  assign s_24 = s_856?s_25:s_855;
  assign s_25 = s_26[24:1];
  assign s_26 = s_842?s_27:s_841;
  dq #(25, 1) dq_s_27 (clk, s_27, s_28);
  assign s_28 = s_29 + s_840;
  assign s_29 = s_30;
  assign s_30 = s_31[47:24];
  dq #(48, 1) dq_s_31 (clk, s_31, s_32);
  assign s_32 = s_33 << s_105;
  dq #(48, 2) dq_s_33 (clk, s_33, s_34);
  dq #(48, 1) dq_s_34 (clk, s_34, s_35);
  assign s_35 = s_36 >> s_90;
  assign s_36 = s_37[47:0];
  assign s_37 = {s_38,s_85};
  assign s_38 = s_39[16:0];
  dq #(34, 1) dq_s_39 (clk, s_39, s_40);
  assign s_40 = s_41 + s_68;
  dq #(34, 2) dq_s_41 (clk, s_41, s_42);
  assign s_42 = s_43 * s_56;
  assign s_43 = s_44;
  assign s_44 = s_45[33:17];
  assign s_45 = s_46;
  assign s_46 = {s_47,s_55};
  assign s_47 = s_50?s_48:s_49;
  assign s_48 = 1'd0;
  assign s_49 = 1'd1;
  assign s_50 = s_51 == s_54;
  assign s_51 = s_52 - s_53;
  assign s_52 = s_5[30:23];
  assign s_53 = 7'd127;
  assign s_54 = -8'd127;
  assign s_55 = s_5[22:0];
  assign s_56 = s_57[33:17];
  assign s_57 = s_58;
  assign s_58 = {s_59,s_67};
  assign s_59 = s_62?s_60:s_61;
  assign s_60 = 1'd0;
  assign s_61 = 1'd1;
  assign s_62 = s_63 == s_66;
  assign s_63 = s_64 - s_65;
  assign s_64 = s_7[30:23];
  assign s_65 = 7'd127;
  assign s_66 = -8'd127;
  assign s_67 = s_7[22:0];
  assign s_68 = s_69 >> s_84;
  dq #(34, 1) dq_s_69 (clk, s_69, s_70);
  assign s_70 = s_71 + s_75;
  dq #(34, 1) dq_s_71 (clk, s_71, s_72);
  assign s_72 = s_73 * s_74;
  assign s_73 = s_44;
  assign s_74 = s_57[16:0];
  dq #(34, 1) dq_s_75 (clk, s_75, s_76);
  assign s_76 = s_77 + s_80;
  assign s_77 = s_78 * s_56;
  assign s_78 = s_79;
  assign s_79 = s_45[16:0];
  assign s_80 = s_81 >> s_83;
  assign s_81 = s_82 * s_74;
  assign s_82 = s_79;
  assign s_83 = 5'd17;
  assign s_84 = 5'd17;
  dq #(34, 1) dq_s_85 (clk, s_85, s_86);
  assign s_86 = {s_87,s_88};
  assign s_87 = s_69[16:0];
  dq #(17, 2) dq_s_88 (clk, s_88, s_89);
  assign s_89 = s_81[16:0];
  dq #(10, 3) dq_s_90 (clk, s_90, s_91);
  assign s_91 = s_104?s_92:s_93;
  assign s_92 = 1'd0;
  assign s_93 = s_94 - s_95;
  assign s_94 = -10'd126;
  assign s_95 = s_96 + s_103;
  assign s_96 = s_97 + s_100;
  assign s_97 = $signed(s_98);
  assign s_98 = s_50?s_99:s_51;
  assign s_99 = -8'd126;
  assign s_100 = $signed(s_101);
  assign s_101 = s_62?s_102:s_63;
  assign s_102 = -8'd126;
  assign s_103 = 1'd1;
  assign s_104 = s_93[9];
  dq #(10, 1) dq_s_105 (clk, s_105, s_106);
  assign s_106 = s_837?s_107:s_832;
  dq #(7, 1) dq_s_107 (clk, s_107, s_108);
  assign s_108 = {s_109,s_826};
  assign s_109 = s_110 & s_484;
  assign s_110 = s_111[5];
  assign s_111 = {s_112,s_478};
  assign s_112 = s_113 & s_312;
  assign s_113 = s_114[4];
  assign s_114 = {s_115,s_306};
  assign s_115 = s_116 & s_228;
  assign s_116 = s_117[3];
  assign s_117 = {s_118,s_222};
  assign s_118 = s_119 & s_188;
  assign s_119 = s_120[2];
  assign s_120 = {s_121,s_182};
  assign s_121 = s_122 & s_170;
  assign s_122 = s_123[1];
  assign s_123 = {s_124,s_166};
  assign s_124 = s_125 & s_164;
  assign s_125 = ~s_126;
  assign s_126 = s_127[1];
  assign s_127 = s_128[3:2];
  assign s_128 = s_129[7:4];
  assign s_129 = s_130[15:8];
  assign s_130 = s_131[31:16];
  assign s_131 = s_132[63:32];
  assign s_132 = {s_133,s_163};
  assign s_133 = {s_134,s_162};
  assign s_134 = {s_135,s_161};
  assign s_135 = {s_136,s_160};
  assign s_136 = {s_137,s_159};
  assign s_137 = {s_138,s_158};
  assign s_138 = {s_139,s_157};
  assign s_139 = {s_140,s_156};
  assign s_140 = {s_141,s_155};
  assign s_141 = {s_142,s_154};
  assign s_142 = {s_143,s_153};
  assign s_143 = {s_144,s_152};
  assign s_144 = {s_145,s_151};
  assign s_145 = {s_146,s_150};
  assign s_146 = {s_147,s_149};
  assign s_147 = {s_34,s_148};
  assign s_148 = 1'd1;
  assign s_149 = 1'd1;
  assign s_150 = 1'd1;
  assign s_151 = 1'd1;
  assign s_152 = 1'd1;
  assign s_153 = 1'd1;
  assign s_154 = 1'd1;
  assign s_155 = 1'd1;
  assign s_156 = 1'd1;
  assign s_157 = 1'd1;
  assign s_158 = 1'd1;
  assign s_159 = 1'd1;
  assign s_160 = 1'd1;
  assign s_161 = 1'd1;
  assign s_162 = 1'd1;
  assign s_163 = 1'd1;
  assign s_164 = ~s_165;
  assign s_165 = s_127[0];
  assign s_166 = s_167 & s_169;
  assign s_167 = ~s_168;
  assign s_168 = s_127[1];
  assign s_169 = s_127[0];
  assign s_170 = s_171[1];
  assign s_171 = {s_172,s_178};
  assign s_172 = s_173 & s_176;
  assign s_173 = ~s_174;
  assign s_174 = s_175[1];
  assign s_175 = s_128[1:0];
  assign s_176 = ~s_177;
  assign s_177 = s_175[0];
  assign s_178 = s_179 & s_181;
  assign s_179 = ~s_180;
  assign s_180 = s_175[1];
  assign s_181 = s_175[0];
  assign s_182 = {s_183,s_185};
  assign s_183 = s_122 & s_184;
  assign s_184 = ~s_170;
  assign s_185 = s_122?s_186:s_187;
  assign s_186 = s_171[0:0];
  assign s_187 = s_123[0:0];
  assign s_188 = s_189[2];
  assign s_189 = {s_190,s_216};
  assign s_190 = s_191 & s_204;
  assign s_191 = s_192[1];
  assign s_192 = {s_193,s_200};
  assign s_193 = s_194 & s_198;
  assign s_194 = ~s_195;
  assign s_195 = s_196[1];
  assign s_196 = s_197[3:2];
  assign s_197 = s_129[3:0];
  assign s_198 = ~s_199;
  assign s_199 = s_196[0];
  assign s_200 = s_201 & s_203;
  assign s_201 = ~s_202;
  assign s_202 = s_196[1];
  assign s_203 = s_196[0];
  assign s_204 = s_205[1];
  assign s_205 = {s_206,s_212};
  assign s_206 = s_207 & s_210;
  assign s_207 = ~s_208;
  assign s_208 = s_209[1];
  assign s_209 = s_197[1:0];
  assign s_210 = ~s_211;
  assign s_211 = s_209[0];
  assign s_212 = s_213 & s_215;
  assign s_213 = ~s_214;
  assign s_214 = s_209[1];
  assign s_215 = s_209[0];
  assign s_216 = {s_217,s_219};
  assign s_217 = s_191 & s_218;
  assign s_218 = ~s_204;
  assign s_219 = s_191?s_220:s_221;
  assign s_220 = s_205[0:0];
  assign s_221 = s_192[0:0];
  assign s_222 = {s_223,s_225};
  assign s_223 = s_119 & s_224;
  assign s_224 = ~s_188;
  assign s_225 = s_119?s_226:s_227;
  assign s_226 = s_189[1:0];
  assign s_227 = s_120[1:0];
  assign s_228 = s_229[3];
  assign s_229 = {s_230,s_300};
  assign s_230 = s_231 & s_266;
  assign s_231 = s_232[2];
  assign s_232 = {s_233,s_260};
  assign s_233 = s_234 & s_248;
  assign s_234 = s_235[1];
  assign s_235 = {s_236,s_244};
  assign s_236 = s_237 & s_242;
  assign s_237 = ~s_238;
  assign s_238 = s_239[1];
  assign s_239 = s_240[3:2];
  assign s_240 = s_241[7:4];
  assign s_241 = s_130[7:0];
  assign s_242 = ~s_243;
  assign s_243 = s_239[0];
  assign s_244 = s_245 & s_247;
  assign s_245 = ~s_246;
  assign s_246 = s_239[1];
  assign s_247 = s_239[0];
  assign s_248 = s_249[1];
  assign s_249 = {s_250,s_256};
  assign s_250 = s_251 & s_254;
  assign s_251 = ~s_252;
  assign s_252 = s_253[1];
  assign s_253 = s_240[1:0];
  assign s_254 = ~s_255;
  assign s_255 = s_253[0];
  assign s_256 = s_257 & s_259;
  assign s_257 = ~s_258;
  assign s_258 = s_253[1];
  assign s_259 = s_253[0];
  assign s_260 = {s_261,s_263};
  assign s_261 = s_234 & s_262;
  assign s_262 = ~s_248;
  assign s_263 = s_234?s_264:s_265;
  assign s_264 = s_249[0:0];
  assign s_265 = s_235[0:0];
  assign s_266 = s_267[2];
  assign s_267 = {s_268,s_294};
  assign s_268 = s_269 & s_282;
  assign s_269 = s_270[1];
  assign s_270 = {s_271,s_278};
  assign s_271 = s_272 & s_276;
  assign s_272 = ~s_273;
  assign s_273 = s_274[1];
  assign s_274 = s_275[3:2];
  assign s_275 = s_241[3:0];
  assign s_276 = ~s_277;
  assign s_277 = s_274[0];
  assign s_278 = s_279 & s_281;
  assign s_279 = ~s_280;
  assign s_280 = s_274[1];
  assign s_281 = s_274[0];
  assign s_282 = s_283[1];
  assign s_283 = {s_284,s_290};
  assign s_284 = s_285 & s_288;
  assign s_285 = ~s_286;
  assign s_286 = s_287[1];
  assign s_287 = s_275[1:0];
  assign s_288 = ~s_289;
  assign s_289 = s_287[0];
  assign s_290 = s_291 & s_293;
  assign s_291 = ~s_292;
  assign s_292 = s_287[1];
  assign s_293 = s_287[0];
  assign s_294 = {s_295,s_297};
  assign s_295 = s_269 & s_296;
  assign s_296 = ~s_282;
  assign s_297 = s_269?s_298:s_299;
  assign s_298 = s_283[0:0];
  assign s_299 = s_270[0:0];
  assign s_300 = {s_301,s_303};
  assign s_301 = s_231 & s_302;
  assign s_302 = ~s_266;
  assign s_303 = s_231?s_304:s_305;
  assign s_304 = s_267[1:0];
  assign s_305 = s_232[1:0];
  assign s_306 = {s_307,s_309};
  assign s_307 = s_116 & s_308;
  assign s_308 = ~s_228;
  assign s_309 = s_116?s_310:s_311;
  assign s_310 = s_229[2:0];
  assign s_311 = s_117[2:0];
  assign s_312 = s_313[4];
  assign s_313 = {s_314,s_472};
  assign s_314 = s_315 & s_394;
  assign s_315 = s_316[3];
  assign s_316 = {s_317,s_388};
  assign s_317 = s_318 & s_354;
  assign s_318 = s_319[2];
  assign s_319 = {s_320,s_348};
  assign s_320 = s_321 & s_336;
  assign s_321 = s_322[1];
  assign s_322 = {s_323,s_332};
  assign s_323 = s_324 & s_330;
  assign s_324 = ~s_325;
  assign s_325 = s_326[1];
  assign s_326 = s_327[3:2];
  assign s_327 = s_328[7:4];
  assign s_328 = s_329[15:8];
  assign s_329 = s_131[15:0];
  assign s_330 = ~s_331;
  assign s_331 = s_326[0];
  assign s_332 = s_333 & s_335;
  assign s_333 = ~s_334;
  assign s_334 = s_326[1];
  assign s_335 = s_326[0];
  assign s_336 = s_337[1];
  assign s_337 = {s_338,s_344};
  assign s_338 = s_339 & s_342;
  assign s_339 = ~s_340;
  assign s_340 = s_341[1];
  assign s_341 = s_327[1:0];
  assign s_342 = ~s_343;
  assign s_343 = s_341[0];
  assign s_344 = s_345 & s_347;
  assign s_345 = ~s_346;
  assign s_346 = s_341[1];
  assign s_347 = s_341[0];
  assign s_348 = {s_349,s_351};
  assign s_349 = s_321 & s_350;
  assign s_350 = ~s_336;
  assign s_351 = s_321?s_352:s_353;
  assign s_352 = s_337[0:0];
  assign s_353 = s_322[0:0];
  assign s_354 = s_355[2];
  assign s_355 = {s_356,s_382};
  assign s_356 = s_357 & s_370;
  assign s_357 = s_358[1];
  assign s_358 = {s_359,s_366};
  assign s_359 = s_360 & s_364;
  assign s_360 = ~s_361;
  assign s_361 = s_362[1];
  assign s_362 = s_363[3:2];
  assign s_363 = s_328[3:0];
  assign s_364 = ~s_365;
  assign s_365 = s_362[0];
  assign s_366 = s_367 & s_369;
  assign s_367 = ~s_368;
  assign s_368 = s_362[1];
  assign s_369 = s_362[0];
  assign s_370 = s_371[1];
  assign s_371 = {s_372,s_378};
  assign s_372 = s_373 & s_376;
  assign s_373 = ~s_374;
  assign s_374 = s_375[1];
  assign s_375 = s_363[1:0];
  assign s_376 = ~s_377;
  assign s_377 = s_375[0];
  assign s_378 = s_379 & s_381;
  assign s_379 = ~s_380;
  assign s_380 = s_375[1];
  assign s_381 = s_375[0];
  assign s_382 = {s_383,s_385};
  assign s_383 = s_357 & s_384;
  assign s_384 = ~s_370;
  assign s_385 = s_357?s_386:s_387;
  assign s_386 = s_371[0:0];
  assign s_387 = s_358[0:0];
  assign s_388 = {s_389,s_391};
  assign s_389 = s_318 & s_390;
  assign s_390 = ~s_354;
  assign s_391 = s_318?s_392:s_393;
  assign s_392 = s_355[1:0];
  assign s_393 = s_319[1:0];
  assign s_394 = s_395[3];
  assign s_395 = {s_396,s_466};
  assign s_396 = s_397 & s_432;
  assign s_397 = s_398[2];
  assign s_398 = {s_399,s_426};
  assign s_399 = s_400 & s_414;
  assign s_400 = s_401[1];
  assign s_401 = {s_402,s_410};
  assign s_402 = s_403 & s_408;
  assign s_403 = ~s_404;
  assign s_404 = s_405[1];
  assign s_405 = s_406[3:2];
  assign s_406 = s_407[7:4];
  assign s_407 = s_329[7:0];
  assign s_408 = ~s_409;
  assign s_409 = s_405[0];
  assign s_410 = s_411 & s_413;
  assign s_411 = ~s_412;
  assign s_412 = s_405[1];
  assign s_413 = s_405[0];
  assign s_414 = s_415[1];
  assign s_415 = {s_416,s_422};
  assign s_416 = s_417 & s_420;
  assign s_417 = ~s_418;
  assign s_418 = s_419[1];
  assign s_419 = s_406[1:0];
  assign s_420 = ~s_421;
  assign s_421 = s_419[0];
  assign s_422 = s_423 & s_425;
  assign s_423 = ~s_424;
  assign s_424 = s_419[1];
  assign s_425 = s_419[0];
  assign s_426 = {s_427,s_429};
  assign s_427 = s_400 & s_428;
  assign s_428 = ~s_414;
  assign s_429 = s_400?s_430:s_431;
  assign s_430 = s_415[0:0];
  assign s_431 = s_401[0:0];
  assign s_432 = s_433[2];
  assign s_433 = {s_434,s_460};
  assign s_434 = s_435 & s_448;
  assign s_435 = s_436[1];
  assign s_436 = {s_437,s_444};
  assign s_437 = s_438 & s_442;
  assign s_438 = ~s_439;
  assign s_439 = s_440[1];
  assign s_440 = s_441[3:2];
  assign s_441 = s_407[3:0];
  assign s_442 = ~s_443;
  assign s_443 = s_440[0];
  assign s_444 = s_445 & s_447;
  assign s_445 = ~s_446;
  assign s_446 = s_440[1];
  assign s_447 = s_440[0];
  assign s_448 = s_449[1];
  assign s_449 = {s_450,s_456};
  assign s_450 = s_451 & s_454;
  assign s_451 = ~s_452;
  assign s_452 = s_453[1];
  assign s_453 = s_441[1:0];
  assign s_454 = ~s_455;
  assign s_455 = s_453[0];
  assign s_456 = s_457 & s_459;
  assign s_457 = ~s_458;
  assign s_458 = s_453[1];
  assign s_459 = s_453[0];
  assign s_460 = {s_461,s_463};
  assign s_461 = s_435 & s_462;
  assign s_462 = ~s_448;
  assign s_463 = s_435?s_464:s_465;
  assign s_464 = s_449[0:0];
  assign s_465 = s_436[0:0];
  assign s_466 = {s_467,s_469};
  assign s_467 = s_397 & s_468;
  assign s_468 = ~s_432;
  assign s_469 = s_397?s_470:s_471;
  assign s_470 = s_433[1:0];
  assign s_471 = s_398[1:0];
  assign s_472 = {s_473,s_475};
  assign s_473 = s_315 & s_474;
  assign s_474 = ~s_394;
  assign s_475 = s_315?s_476:s_477;
  assign s_476 = s_395[2:0];
  assign s_477 = s_316[2:0];
  assign s_478 = {s_479,s_481};
  assign s_479 = s_113 & s_480;
  assign s_480 = ~s_312;
  assign s_481 = s_113?s_482:s_483;
  assign s_482 = s_313[3:0];
  assign s_483 = s_114[3:0];
  assign s_484 = s_485[5];
  assign s_485 = {s_486,s_820};
  assign s_486 = s_487 & s_654;
  assign s_487 = s_488[4];
  assign s_488 = {s_489,s_648};
  assign s_489 = s_490 & s_570;
  assign s_490 = s_491[3];
  assign s_491 = {s_492,s_564};
  assign s_492 = s_493 & s_530;
  assign s_493 = s_494[2];
  assign s_494 = {s_495,s_524};
  assign s_495 = s_496 & s_512;
  assign s_496 = s_497[1];
  assign s_497 = {s_498,s_508};
  assign s_498 = s_499 & s_506;
  assign s_499 = ~s_500;
  assign s_500 = s_501[1];
  assign s_501 = s_502[3:2];
  assign s_502 = s_503[7:4];
  assign s_503 = s_504[15:8];
  assign s_504 = s_505[31:16];
  assign s_505 = s_132[31:0];
  assign s_506 = ~s_507;
  assign s_507 = s_501[0];
  assign s_508 = s_509 & s_511;
  assign s_509 = ~s_510;
  assign s_510 = s_501[1];
  assign s_511 = s_501[0];
  assign s_512 = s_513[1];
  assign s_513 = {s_514,s_520};
  assign s_514 = s_515 & s_518;
  assign s_515 = ~s_516;
  assign s_516 = s_517[1];
  assign s_517 = s_502[1:0];
  assign s_518 = ~s_519;
  assign s_519 = s_517[0];
  assign s_520 = s_521 & s_523;
  assign s_521 = ~s_522;
  assign s_522 = s_517[1];
  assign s_523 = s_517[0];
  assign s_524 = {s_525,s_527};
  assign s_525 = s_496 & s_526;
  assign s_526 = ~s_512;
  assign s_527 = s_496?s_528:s_529;
  assign s_528 = s_513[0:0];
  assign s_529 = s_497[0:0];
  assign s_530 = s_531[2];
  assign s_531 = {s_532,s_558};
  assign s_532 = s_533 & s_546;
  assign s_533 = s_534[1];
  assign s_534 = {s_535,s_542};
  assign s_535 = s_536 & s_540;
  assign s_536 = ~s_537;
  assign s_537 = s_538[1];
  assign s_538 = s_539[3:2];
  assign s_539 = s_503[3:0];
  assign s_540 = ~s_541;
  assign s_541 = s_538[0];
  assign s_542 = s_543 & s_545;
  assign s_543 = ~s_544;
  assign s_544 = s_538[1];
  assign s_545 = s_538[0];
  assign s_546 = s_547[1];
  assign s_547 = {s_548,s_554};
  assign s_548 = s_549 & s_552;
  assign s_549 = ~s_550;
  assign s_550 = s_551[1];
  assign s_551 = s_539[1:0];
  assign s_552 = ~s_553;
  assign s_553 = s_551[0];
  assign s_554 = s_555 & s_557;
  assign s_555 = ~s_556;
  assign s_556 = s_551[1];
  assign s_557 = s_551[0];
  assign s_558 = {s_559,s_561};
  assign s_559 = s_533 & s_560;
  assign s_560 = ~s_546;
  assign s_561 = s_533?s_562:s_563;
  assign s_562 = s_547[0:0];
  assign s_563 = s_534[0:0];
  assign s_564 = {s_565,s_567};
  assign s_565 = s_493 & s_566;
  assign s_566 = ~s_530;
  assign s_567 = s_493?s_568:s_569;
  assign s_568 = s_531[1:0];
  assign s_569 = s_494[1:0];
  assign s_570 = s_571[3];
  assign s_571 = {s_572,s_642};
  assign s_572 = s_573 & s_608;
  assign s_573 = s_574[2];
  assign s_574 = {s_575,s_602};
  assign s_575 = s_576 & s_590;
  assign s_576 = s_577[1];
  assign s_577 = {s_578,s_586};
  assign s_578 = s_579 & s_584;
  assign s_579 = ~s_580;
  assign s_580 = s_581[1];
  assign s_581 = s_582[3:2];
  assign s_582 = s_583[7:4];
  assign s_583 = s_504[7:0];
  assign s_584 = ~s_585;
  assign s_585 = s_581[0];
  assign s_586 = s_587 & s_589;
  assign s_587 = ~s_588;
  assign s_588 = s_581[1];
  assign s_589 = s_581[0];
  assign s_590 = s_591[1];
  assign s_591 = {s_592,s_598};
  assign s_592 = s_593 & s_596;
  assign s_593 = ~s_594;
  assign s_594 = s_595[1];
  assign s_595 = s_582[1:0];
  assign s_596 = ~s_597;
  assign s_597 = s_595[0];
  assign s_598 = s_599 & s_601;
  assign s_599 = ~s_600;
  assign s_600 = s_595[1];
  assign s_601 = s_595[0];
  assign s_602 = {s_603,s_605};
  assign s_603 = s_576 & s_604;
  assign s_604 = ~s_590;
  assign s_605 = s_576?s_606:s_607;
  assign s_606 = s_591[0:0];
  assign s_607 = s_577[0:0];
  assign s_608 = s_609[2];
  assign s_609 = {s_610,s_636};
  assign s_610 = s_611 & s_624;
  assign s_611 = s_612[1];
  assign s_612 = {s_613,s_620};
  assign s_613 = s_614 & s_618;
  assign s_614 = ~s_615;
  assign s_615 = s_616[1];
  assign s_616 = s_617[3:2];
  assign s_617 = s_583[3:0];
  assign s_618 = ~s_619;
  assign s_619 = s_616[0];
  assign s_620 = s_621 & s_623;
  assign s_621 = ~s_622;
  assign s_622 = s_616[1];
  assign s_623 = s_616[0];
  assign s_624 = s_625[1];
  assign s_625 = {s_626,s_632};
  assign s_626 = s_627 & s_630;
  assign s_627 = ~s_628;
  assign s_628 = s_629[1];
  assign s_629 = s_617[1:0];
  assign s_630 = ~s_631;
  assign s_631 = s_629[0];
  assign s_632 = s_633 & s_635;
  assign s_633 = ~s_634;
  assign s_634 = s_629[1];
  assign s_635 = s_629[0];
  assign s_636 = {s_637,s_639};
  assign s_637 = s_611 & s_638;
  assign s_638 = ~s_624;
  assign s_639 = s_611?s_640:s_641;
  assign s_640 = s_625[0:0];
  assign s_641 = s_612[0:0];
  assign s_642 = {s_643,s_645};
  assign s_643 = s_573 & s_644;
  assign s_644 = ~s_608;
  assign s_645 = s_573?s_646:s_647;
  assign s_646 = s_609[1:0];
  assign s_647 = s_574[1:0];
  assign s_648 = {s_649,s_651};
  assign s_649 = s_490 & s_650;
  assign s_650 = ~s_570;
  assign s_651 = s_490?s_652:s_653;
  assign s_652 = s_571[2:0];
  assign s_653 = s_491[2:0];
  assign s_654 = s_655[4];
  assign s_655 = {s_656,s_814};
  assign s_656 = s_657 & s_736;
  assign s_657 = s_658[3];
  assign s_658 = {s_659,s_730};
  assign s_659 = s_660 & s_696;
  assign s_660 = s_661[2];
  assign s_661 = {s_662,s_690};
  assign s_662 = s_663 & s_678;
  assign s_663 = s_664[1];
  assign s_664 = {s_665,s_674};
  assign s_665 = s_666 & s_672;
  assign s_666 = ~s_667;
  assign s_667 = s_668[1];
  assign s_668 = s_669[3:2];
  assign s_669 = s_670[7:4];
  assign s_670 = s_671[15:8];
  assign s_671 = s_505[15:0];
  assign s_672 = ~s_673;
  assign s_673 = s_668[0];
  assign s_674 = s_675 & s_677;
  assign s_675 = ~s_676;
  assign s_676 = s_668[1];
  assign s_677 = s_668[0];
  assign s_678 = s_679[1];
  assign s_679 = {s_680,s_686};
  assign s_680 = s_681 & s_684;
  assign s_681 = ~s_682;
  assign s_682 = s_683[1];
  assign s_683 = s_669[1:0];
  assign s_684 = ~s_685;
  assign s_685 = s_683[0];
  assign s_686 = s_687 & s_689;
  assign s_687 = ~s_688;
  assign s_688 = s_683[1];
  assign s_689 = s_683[0];
  assign s_690 = {s_691,s_693};
  assign s_691 = s_663 & s_692;
  assign s_692 = ~s_678;
  assign s_693 = s_663?s_694:s_695;
  assign s_694 = s_679[0:0];
  assign s_695 = s_664[0:0];
  assign s_696 = s_697[2];
  assign s_697 = {s_698,s_724};
  assign s_698 = s_699 & s_712;
  assign s_699 = s_700[1];
  assign s_700 = {s_701,s_708};
  assign s_701 = s_702 & s_706;
  assign s_702 = ~s_703;
  assign s_703 = s_704[1];
  assign s_704 = s_705[3:2];
  assign s_705 = s_670[3:0];
  assign s_706 = ~s_707;
  assign s_707 = s_704[0];
  assign s_708 = s_709 & s_711;
  assign s_709 = ~s_710;
  assign s_710 = s_704[1];
  assign s_711 = s_704[0];
  assign s_712 = s_713[1];
  assign s_713 = {s_714,s_720};
  assign s_714 = s_715 & s_718;
  assign s_715 = ~s_716;
  assign s_716 = s_717[1];
  assign s_717 = s_705[1:0];
  assign s_718 = ~s_719;
  assign s_719 = s_717[0];
  assign s_720 = s_721 & s_723;
  assign s_721 = ~s_722;
  assign s_722 = s_717[1];
  assign s_723 = s_717[0];
  assign s_724 = {s_725,s_727};
  assign s_725 = s_699 & s_726;
  assign s_726 = ~s_712;
  assign s_727 = s_699?s_728:s_729;
  assign s_728 = s_713[0:0];
  assign s_729 = s_700[0:0];
  assign s_730 = {s_731,s_733};
  assign s_731 = s_660 & s_732;
  assign s_732 = ~s_696;
  assign s_733 = s_660?s_734:s_735;
  assign s_734 = s_697[1:0];
  assign s_735 = s_661[1:0];
  assign s_736 = s_737[3];
  assign s_737 = {s_738,s_808};
  assign s_738 = s_739 & s_774;
  assign s_739 = s_740[2];
  assign s_740 = {s_741,s_768};
  assign s_741 = s_742 & s_756;
  assign s_742 = s_743[1];
  assign s_743 = {s_744,s_752};
  assign s_744 = s_745 & s_750;
  assign s_745 = ~s_746;
  assign s_746 = s_747[1];
  assign s_747 = s_748[3:2];
  assign s_748 = s_749[7:4];
  assign s_749 = s_671[7:0];
  assign s_750 = ~s_751;
  assign s_751 = s_747[0];
  assign s_752 = s_753 & s_755;
  assign s_753 = ~s_754;
  assign s_754 = s_747[1];
  assign s_755 = s_747[0];
  assign s_756 = s_757[1];
  assign s_757 = {s_758,s_764};
  assign s_758 = s_759 & s_762;
  assign s_759 = ~s_760;
  assign s_760 = s_761[1];
  assign s_761 = s_748[1:0];
  assign s_762 = ~s_763;
  assign s_763 = s_761[0];
  assign s_764 = s_765 & s_767;
  assign s_765 = ~s_766;
  assign s_766 = s_761[1];
  assign s_767 = s_761[0];
  assign s_768 = {s_769,s_771};
  assign s_769 = s_742 & s_770;
  assign s_770 = ~s_756;
  assign s_771 = s_742?s_772:s_773;
  assign s_772 = s_757[0:0];
  assign s_773 = s_743[0:0];
  assign s_774 = s_775[2];
  assign s_775 = {s_776,s_802};
  assign s_776 = s_777 & s_790;
  assign s_777 = s_778[1];
  assign s_778 = {s_779,s_786};
  assign s_779 = s_780 & s_784;
  assign s_780 = ~s_781;
  assign s_781 = s_782[1];
  assign s_782 = s_783[3:2];
  assign s_783 = s_749[3:0];
  assign s_784 = ~s_785;
  assign s_785 = s_782[0];
  assign s_786 = s_787 & s_789;
  assign s_787 = ~s_788;
  assign s_788 = s_782[1];
  assign s_789 = s_782[0];
  assign s_790 = s_791[1];
  assign s_791 = {s_792,s_798};
  assign s_792 = s_793 & s_796;
  assign s_793 = ~s_794;
  assign s_794 = s_795[1];
  assign s_795 = s_783[1:0];
  assign s_796 = ~s_797;
  assign s_797 = s_795[0];
  assign s_798 = s_799 & s_801;
  assign s_799 = ~s_800;
  assign s_800 = s_795[1];
  assign s_801 = s_795[0];
  assign s_802 = {s_803,s_805};
  assign s_803 = s_777 & s_804;
  assign s_804 = ~s_790;
  assign s_805 = s_777?s_806:s_807;
  assign s_806 = s_791[0:0];
  assign s_807 = s_778[0:0];
  assign s_808 = {s_809,s_811};
  assign s_809 = s_739 & s_810;
  assign s_810 = ~s_774;
  assign s_811 = s_739?s_812:s_813;
  assign s_812 = s_775[1:0];
  assign s_813 = s_740[1:0];
  assign s_814 = {s_815,s_817};
  assign s_815 = s_657 & s_816;
  assign s_816 = ~s_736;
  assign s_817 = s_657?s_818:s_819;
  assign s_818 = s_737[2:0];
  assign s_819 = s_658[2:0];
  assign s_820 = {s_821,s_823};
  assign s_821 = s_487 & s_822;
  assign s_822 = ~s_654;
  assign s_823 = s_487?s_824:s_825;
  assign s_824 = s_655[3:0];
  assign s_825 = s_488[3:0];
  assign s_826 = {s_827,s_829};
  assign s_827 = s_110 & s_828;
  assign s_828 = ~s_484;
  assign s_829 = s_110?s_830:s_831;
  assign s_830 = s_485[4:0];
  assign s_831 = s_111[4:0];
  dq #(10, 4) dq_s_832 (clk, s_832, s_833);
  assign s_833 = s_834 - s_836;
  dq #(10, 1) dq_s_834 (clk, s_834, s_835);
  assign s_835 = s_95 + s_91;
  assign s_836 = -10'd126;
  assign s_837 = s_838 <= s_839;
  assign s_838 = s_107;
  dq #(10, 4) dq_s_839 (clk, s_839, s_833);
  assign s_840 = 1'd1;
  dq #(24, 1) dq_s_841 (clk, s_841, s_30);
  assign s_842 = s_843 & s_845;
  dq #(1, 1) dq_s_843 (clk, s_843, s_844);
  assign s_844 = s_31[23];
  assign s_845 = s_846 | s_853;
  assign s_846 = s_847 | s_849;
  dq #(1, 1) dq_s_847 (clk, s_847, s_848);
  assign s_848 = s_31[22];
  dq #(1, 1) dq_s_849 (clk, s_849, s_850);
  assign s_850 = s_851 != s_852;
  assign s_851 = s_31[21:0];
  assign s_852 = 24'd0;
  dq #(1, 1) dq_s_853 (clk, s_853, s_854);
  assign s_854 = s_30[0];
  assign s_855 = s_26[23:0];
  assign s_856 = s_26[24];
  assign s_857 = {s_858,s_869};
  assign s_858 = {s_859,s_860};
  dq #(1, 9) dq_s_859 (clk, s_859, s_3);
  assign s_860 = s_861 + s_868;
  assign s_861 = s_862[7:0];
  dq #(10, 1) dq_s_862 (clk, s_862, s_863);
  assign s_863 = s_864 + s_856;
  dq #(10, 1) dq_s_864 (clk, s_864, s_865);
  dq #(10, 1) dq_s_865 (clk, s_865, s_866);
  assign s_866 = s_867 - s_105;
  dq #(10, 5) dq_s_867 (clk, s_867, s_834);
  assign s_868 = 7'd127;
  assign s_869 = s_23[22:0];
  assign s_870 = s_871 & s_873;
  assign s_871 = s_861 == s_872;
  assign s_872 = -8'd126;
  assign s_873 = ~s_874;
  assign s_874 = s_23[23];
  assign s_875 = s_23 == s_876;
  assign s_876 = 24'd0;
  assign s_877 = s_878 | s_887;
  assign s_878 = s_879 | s_881;
  assign s_879 = $signed(s_862) > $signed(s_880);
  assign s_880 = 9'd127;
  dq #(1, 9) dq_s_881 (clk, s_881, s_882);
  assign s_882 = s_883 & s_885;
  assign s_883 = s_51 == s_884;
  assign s_884 = 8'd128;
  assign s_885 = s_55 == s_886;
  assign s_886 = 23'd0;
  dq #(1, 9) dq_s_887 (clk, s_887, s_888);
  assign s_888 = s_889 & s_891;
  assign s_889 = s_63 == s_890;
  assign s_890 = 8'd128;
  assign s_891 = s_67 == s_892;
  assign s_892 = 23'd0;
  dq #(1, 9) dq_s_893 (clk, s_893, s_894);
  assign s_894 = s_895 | s_900;
  assign s_895 = s_896 & s_898;
  assign s_896 = s_51 == s_897;
  assign s_897 = 8'd128;
  assign s_898 = s_55 != s_899;
  assign s_899 = 23'd0;
  assign s_900 = s_901 & s_903;
  assign s_901 = s_63 == s_902;
  assign s_902 = 8'd128;
  assign s_903 = s_67 != s_904;
  assign s_904 = 23'd0;
  assign mul_z = s_0;
endmodule
