module dq (clk, q, d);
  input  clk;
  input  [width-1:0] d;
  output [width-1:0] q;
  parameter width=8;
  parameter depth=2;
  integer i;
  reg [width-1:0] delay_line [depth-1:0];
  always @(posedge clk) begin
    delay_line[0] <= d;
    for(i=1; i<depth; i=i+1) begin
      delay_line[i] <= delay_line[i-1];
    end
  end
  assign q = delay_line[depth-1];
endmodule

module double_sqrt(clk, double_sqrt_a, double_sqrt_z);
  input clk;
  input [63:0] double_sqrt_a;
  output [63:0] double_sqrt_z;
  wire [63:0] s_0;
  wire [63:0] s_1;
  wire [63:0] s_2;
  wire [0:0] s_3;
  wire [63:0] s_4;
  wire [62:0] s_5;
  wire [63:0] s_6;
  wire [63:0] s_7;
  wire [63:0] s_8;
  wire [62:0] s_9;
  wire [63:0] s_10;
  wire [63:0] s_11;
  wire [63:0] s_12;
  wire [62:0] s_13;
  wire [63:0] s_14;
  wire [63:0] s_15;
  wire [11:0] s_16;
  wire [11:0] s_17;
  wire [10:0] s_18;
  wire [51:0] s_19;
  wire [52:0] s_20;
  wire [52:0] s_21;
  wire [52:0] s_22;
  wire [53:0] s_23;
  wire [53:0] s_24;
  wire [53:0] s_25;
  wire [52:0] s_26;
  wire [53:0] s_27;
  wire [53:0] s_28;
  wire [53:0] s_29;
  wire [53:0] s_30;
  wire [53:0] s_31;
  wire [53:0] s_32;
  wire [53:0] s_33;
  wire [108:0] s_34;
  wire [108:0] s_35;
  wire [108:0] s_36;
  wire [108:0] s_37;
  wire [108:0] s_38;
  wire [108:0] s_39;
  wire [108:0] s_40;
  wire [108:0] s_41;
  wire [108:0] s_42;
  wire [108:0] s_43;
  wire [108:0] s_44;
  wire [108:0] s_45;
  wire [108:0] s_46;
  wire [108:0] s_47;
  wire [108:0] s_48;
  wire [108:0] s_49;
  wire [108:0] s_50;
  wire [108:0] s_51;
  wire [108:0] s_52;
  wire [108:0] s_53;
  wire [108:0] s_54;
  wire [108:0] s_55;
  wire [108:0] s_56;
  wire [108:0] s_57;
  wire [108:0] s_58;
  wire [108:0] s_59;
  wire [108:0] s_60;
  wire [108:0] s_61;
  wire [108:0] s_62;
  wire [108:0] s_63;
  wire [108:0] s_64;
  wire [108:0] s_65;
  wire [108:0] s_66;
  wire [108:0] s_67;
  wire [108:0] s_68;
  wire [108:0] s_69;
  wire [108:0] s_70;
  wire [108:0] s_71;
  wire [108:0] s_72;
  wire [108:0] s_73;
  wire [108:0] s_74;
  wire [108:0] s_75;
  wire [108:0] s_76;
  wire [108:0] s_77;
  wire [108:0] s_78;
  wire [108:0] s_79;
  wire [108:0] s_80;
  wire [108:0] s_81;
  wire [108:0] s_82;
  wire [108:0] s_83;
  wire [108:0] s_84;
  wire [108:0] s_85;
  wire [108:0] s_86;
  wire [108:0] s_87;
  wire [108:0] s_88;
  wire [108:0] s_89;
  wire [108:0] s_90;
  wire [108:0] s_91;
  wire [108:0] s_92;
  wire [108:0] s_93;
  wire [108:0] s_94;
  wire [108:0] s_95;
  wire [108:0] s_96;
  wire [108:0] s_97;
  wire [108:0] s_98;
  wire [108:0] s_99;
  wire [108:0] s_100;
  wire [108:0] s_101;
  wire [108:0] s_102;
  wire [108:0] s_103;
  wire [108:0] s_104;
  wire [108:0] s_105;
  wire [108:0] s_106;
  wire [108:0] s_107;
  wire [108:0] s_108;
  wire [108:0] s_109;
  wire [108:0] s_110;
  wire [108:0] s_111;
  wire [108:0] s_112;
  wire [108:0] s_113;
  wire [108:0] s_114;
  wire [108:0] s_115;
  wire [108:0] s_116;
  wire [108:0] s_117;
  wire [108:0] s_118;
  wire [108:0] s_119;
  wire [108:0] s_120;
  wire [108:0] s_121;
  wire [108:0] s_122;
  wire [108:0] s_123;
  wire [108:0] s_124;
  wire [108:0] s_125;
  wire [108:0] s_126;
  wire [108:0] s_127;
  wire [108:0] s_128;
  wire [108:0] s_129;
  wire [108:0] s_130;
  wire [108:0] s_131;
  wire [108:0] s_132;
  wire [108:0] s_133;
  wire [108:0] s_134;
  wire [108:0] s_135;
  wire [108:0] s_136;
  wire [108:0] s_137;
  wire [108:0] s_138;
  wire [108:0] s_139;
  wire [108:0] s_140;
  wire [108:0] s_141;
  wire [108:0] s_142;
  wire [108:0] s_143;
  wire [108:0] s_144;
  wire [54:0] s_145;
  wire [108:0] s_146;
  wire [0:0] s_147;
  wire [109:0] s_148;
  wire [109:0] s_149;
  wire [109:0] s_150;
  wire [109:0] s_151;
  wire [54:0] s_152;
  wire [5:0] s_153;
  wire [108:0] s_154;
  wire [108:0] s_155;
  wire [108:0] s_156;
  wire [108:0] s_157;
  wire [108:0] s_158;
  wire [52:0] s_159;
  wire [52:0] s_160;
  wire [52:0] s_161;
  wire [52:0] s_162;
  wire [0:0] s_163;
  wire [0:0] s_164;
  wire [0:0] s_165;
  wire [0:0] s_166;
  wire [10:0] s_167;
  wire [10:0] s_168;
  wire [9:0] s_169;
  wire [10:0] s_170;
  wire [51:0] s_171;
  wire [12:0] s_172;
  wire [12:0] s_173;
  wire [6:0] s_174;
  wire [6:0] s_175;
  wire [0:0] s_176;
  wire [0:0] s_177;
  wire [5:0] s_178;
  wire [0:0] s_179;
  wire [0:0] s_180;
  wire [4:0] s_181;
  wire [0:0] s_182;
  wire [0:0] s_183;
  wire [3:0] s_184;
  wire [0:0] s_185;
  wire [0:0] s_186;
  wire [2:0] s_187;
  wire [0:0] s_188;
  wire [0:0] s_189;
  wire [1:0] s_190;
  wire [0:0] s_191;
  wire [0:0] s_192;
  wire [0:0] s_193;
  wire [1:0] s_194;
  wire [3:0] s_195;
  wire [7:0] s_196;
  wire [15:0] s_197;
  wire [31:0] s_198;
  wire [63:0] s_199;
  wire [62:0] s_200;
  wire [61:0] s_201;
  wire [60:0] s_202;
  wire [59:0] s_203;
  wire [58:0] s_204;
  wire [57:0] s_205;
  wire [56:0] s_206;
  wire [55:0] s_207;
  wire [54:0] s_208;
  wire [53:0] s_209;
  wire [0:0] s_210;
  wire [0:0] s_211;
  wire [0:0] s_212;
  wire [0:0] s_213;
  wire [0:0] s_214;
  wire [0:0] s_215;
  wire [0:0] s_216;
  wire [0:0] s_217;
  wire [0:0] s_218;
  wire [0:0] s_219;
  wire [0:0] s_220;
  wire [0:0] s_221;
  wire [0:0] s_222;
  wire [0:0] s_223;
  wire [0:0] s_224;
  wire [0:0] s_225;
  wire [0:0] s_226;
  wire [0:0] s_227;
  wire [1:0] s_228;
  wire [0:0] s_229;
  wire [0:0] s_230;
  wire [0:0] s_231;
  wire [1:0] s_232;
  wire [0:0] s_233;
  wire [0:0] s_234;
  wire [0:0] s_235;
  wire [0:0] s_236;
  wire [0:0] s_237;
  wire [0:0] s_238;
  wire [1:0] s_239;
  wire [0:0] s_240;
  wire [0:0] s_241;
  wire [0:0] s_242;
  wire [0:0] s_243;
  wire [0:0] s_244;
  wire [0:0] s_245;
  wire [2:0] s_246;
  wire [0:0] s_247;
  wire [0:0] s_248;
  wire [1:0] s_249;
  wire [0:0] s_250;
  wire [0:0] s_251;
  wire [0:0] s_252;
  wire [1:0] s_253;
  wire [3:0] s_254;
  wire [0:0] s_255;
  wire [0:0] s_256;
  wire [0:0] s_257;
  wire [0:0] s_258;
  wire [0:0] s_259;
  wire [0:0] s_260;
  wire [0:0] s_261;
  wire [1:0] s_262;
  wire [0:0] s_263;
  wire [0:0] s_264;
  wire [0:0] s_265;
  wire [1:0] s_266;
  wire [0:0] s_267;
  wire [0:0] s_268;
  wire [0:0] s_269;
  wire [0:0] s_270;
  wire [0:0] s_271;
  wire [0:0] s_272;
  wire [1:0] s_273;
  wire [0:0] s_274;
  wire [0:0] s_275;
  wire [0:0] s_276;
  wire [0:0] s_277;
  wire [0:0] s_278;
  wire [2:0] s_279;
  wire [0:0] s_280;
  wire [0:0] s_281;
  wire [1:0] s_282;
  wire [1:0] s_283;
  wire [1:0] s_284;
  wire [0:0] s_285;
  wire [3:0] s_286;
  wire [0:0] s_287;
  wire [0:0] s_288;
  wire [2:0] s_289;
  wire [0:0] s_290;
  wire [0:0] s_291;
  wire [1:0] s_292;
  wire [0:0] s_293;
  wire [0:0] s_294;
  wire [0:0] s_295;
  wire [1:0] s_296;
  wire [3:0] s_297;
  wire [7:0] s_298;
  wire [0:0] s_299;
  wire [0:0] s_300;
  wire [0:0] s_301;
  wire [0:0] s_302;
  wire [0:0] s_303;
  wire [0:0] s_304;
  wire [0:0] s_305;
  wire [1:0] s_306;
  wire [0:0] s_307;
  wire [0:0] s_308;
  wire [0:0] s_309;
  wire [1:0] s_310;
  wire [0:0] s_311;
  wire [0:0] s_312;
  wire [0:0] s_313;
  wire [0:0] s_314;
  wire [0:0] s_315;
  wire [0:0] s_316;
  wire [1:0] s_317;
  wire [0:0] s_318;
  wire [0:0] s_319;
  wire [0:0] s_320;
  wire [0:0] s_321;
  wire [0:0] s_322;
  wire [0:0] s_323;
  wire [2:0] s_324;
  wire [0:0] s_325;
  wire [0:0] s_326;
  wire [1:0] s_327;
  wire [0:0] s_328;
  wire [0:0] s_329;
  wire [0:0] s_330;
  wire [1:0] s_331;
  wire [3:0] s_332;
  wire [0:0] s_333;
  wire [0:0] s_334;
  wire [0:0] s_335;
  wire [0:0] s_336;
  wire [0:0] s_337;
  wire [0:0] s_338;
  wire [0:0] s_339;
  wire [1:0] s_340;
  wire [0:0] s_341;
  wire [0:0] s_342;
  wire [0:0] s_343;
  wire [1:0] s_344;
  wire [0:0] s_345;
  wire [0:0] s_346;
  wire [0:0] s_347;
  wire [0:0] s_348;
  wire [0:0] s_349;
  wire [0:0] s_350;
  wire [1:0] s_351;
  wire [0:0] s_352;
  wire [0:0] s_353;
  wire [0:0] s_354;
  wire [0:0] s_355;
  wire [0:0] s_356;
  wire [2:0] s_357;
  wire [0:0] s_358;
  wire [0:0] s_359;
  wire [1:0] s_360;
  wire [1:0] s_361;
  wire [1:0] s_362;
  wire [3:0] s_363;
  wire [0:0] s_364;
  wire [0:0] s_365;
  wire [2:0] s_366;
  wire [2:0] s_367;
  wire [2:0] s_368;
  wire [0:0] s_369;
  wire [4:0] s_370;
  wire [0:0] s_371;
  wire [0:0] s_372;
  wire [3:0] s_373;
  wire [0:0] s_374;
  wire [0:0] s_375;
  wire [2:0] s_376;
  wire [0:0] s_377;
  wire [0:0] s_378;
  wire [1:0] s_379;
  wire [0:0] s_380;
  wire [0:0] s_381;
  wire [0:0] s_382;
  wire [1:0] s_383;
  wire [3:0] s_384;
  wire [7:0] s_385;
  wire [15:0] s_386;
  wire [0:0] s_387;
  wire [0:0] s_388;
  wire [0:0] s_389;
  wire [0:0] s_390;
  wire [0:0] s_391;
  wire [0:0] s_392;
  wire [0:0] s_393;
  wire [1:0] s_394;
  wire [0:0] s_395;
  wire [0:0] s_396;
  wire [0:0] s_397;
  wire [1:0] s_398;
  wire [0:0] s_399;
  wire [0:0] s_400;
  wire [0:0] s_401;
  wire [0:0] s_402;
  wire [0:0] s_403;
  wire [0:0] s_404;
  wire [1:0] s_405;
  wire [0:0] s_406;
  wire [0:0] s_407;
  wire [0:0] s_408;
  wire [0:0] s_409;
  wire [0:0] s_410;
  wire [0:0] s_411;
  wire [2:0] s_412;
  wire [0:0] s_413;
  wire [0:0] s_414;
  wire [1:0] s_415;
  wire [0:0] s_416;
  wire [0:0] s_417;
  wire [0:0] s_418;
  wire [1:0] s_419;
  wire [3:0] s_420;
  wire [0:0] s_421;
  wire [0:0] s_422;
  wire [0:0] s_423;
  wire [0:0] s_424;
  wire [0:0] s_425;
  wire [0:0] s_426;
  wire [0:0] s_427;
  wire [1:0] s_428;
  wire [0:0] s_429;
  wire [0:0] s_430;
  wire [0:0] s_431;
  wire [1:0] s_432;
  wire [0:0] s_433;
  wire [0:0] s_434;
  wire [0:0] s_435;
  wire [0:0] s_436;
  wire [0:0] s_437;
  wire [0:0] s_438;
  wire [1:0] s_439;
  wire [0:0] s_440;
  wire [0:0] s_441;
  wire [0:0] s_442;
  wire [0:0] s_443;
  wire [0:0] s_444;
  wire [2:0] s_445;
  wire [0:0] s_446;
  wire [0:0] s_447;
  wire [1:0] s_448;
  wire [1:0] s_449;
  wire [1:0] s_450;
  wire [0:0] s_451;
  wire [3:0] s_452;
  wire [0:0] s_453;
  wire [0:0] s_454;
  wire [2:0] s_455;
  wire [0:0] s_456;
  wire [0:0] s_457;
  wire [1:0] s_458;
  wire [0:0] s_459;
  wire [0:0] s_460;
  wire [0:0] s_461;
  wire [1:0] s_462;
  wire [3:0] s_463;
  wire [7:0] s_464;
  wire [0:0] s_465;
  wire [0:0] s_466;
  wire [0:0] s_467;
  wire [0:0] s_468;
  wire [0:0] s_469;
  wire [0:0] s_470;
  wire [0:0] s_471;
  wire [1:0] s_472;
  wire [0:0] s_473;
  wire [0:0] s_474;
  wire [0:0] s_475;
  wire [1:0] s_476;
  wire [0:0] s_477;
  wire [0:0] s_478;
  wire [0:0] s_479;
  wire [0:0] s_480;
  wire [0:0] s_481;
  wire [0:0] s_482;
  wire [1:0] s_483;
  wire [0:0] s_484;
  wire [0:0] s_485;
  wire [0:0] s_486;
  wire [0:0] s_487;
  wire [0:0] s_488;
  wire [0:0] s_489;
  wire [2:0] s_490;
  wire [0:0] s_491;
  wire [0:0] s_492;
  wire [1:0] s_493;
  wire [0:0] s_494;
  wire [0:0] s_495;
  wire [0:0] s_496;
  wire [1:0] s_497;
  wire [3:0] s_498;
  wire [0:0] s_499;
  wire [0:0] s_500;
  wire [0:0] s_501;
  wire [0:0] s_502;
  wire [0:0] s_503;
  wire [0:0] s_504;
  wire [0:0] s_505;
  wire [1:0] s_506;
  wire [0:0] s_507;
  wire [0:0] s_508;
  wire [0:0] s_509;
  wire [1:0] s_510;
  wire [0:0] s_511;
  wire [0:0] s_512;
  wire [0:0] s_513;
  wire [0:0] s_514;
  wire [0:0] s_515;
  wire [0:0] s_516;
  wire [1:0] s_517;
  wire [0:0] s_518;
  wire [0:0] s_519;
  wire [0:0] s_520;
  wire [0:0] s_521;
  wire [0:0] s_522;
  wire [2:0] s_523;
  wire [0:0] s_524;
  wire [0:0] s_525;
  wire [1:0] s_526;
  wire [1:0] s_527;
  wire [1:0] s_528;
  wire [3:0] s_529;
  wire [0:0] s_530;
  wire [0:0] s_531;
  wire [2:0] s_532;
  wire [2:0] s_533;
  wire [2:0] s_534;
  wire [4:0] s_535;
  wire [0:0] s_536;
  wire [0:0] s_537;
  wire [3:0] s_538;
  wire [3:0] s_539;
  wire [3:0] s_540;
  wire [0:0] s_541;
  wire [5:0] s_542;
  wire [0:0] s_543;
  wire [0:0] s_544;
  wire [4:0] s_545;
  wire [0:0] s_546;
  wire [0:0] s_547;
  wire [3:0] s_548;
  wire [0:0] s_549;
  wire [0:0] s_550;
  wire [2:0] s_551;
  wire [0:0] s_552;
  wire [0:0] s_553;
  wire [1:0] s_554;
  wire [0:0] s_555;
  wire [0:0] s_556;
  wire [0:0] s_557;
  wire [1:0] s_558;
  wire [3:0] s_559;
  wire [7:0] s_560;
  wire [15:0] s_561;
  wire [31:0] s_562;
  wire [0:0] s_563;
  wire [0:0] s_564;
  wire [0:0] s_565;
  wire [0:0] s_566;
  wire [0:0] s_567;
  wire [0:0] s_568;
  wire [0:0] s_569;
  wire [1:0] s_570;
  wire [0:0] s_571;
  wire [0:0] s_572;
  wire [0:0] s_573;
  wire [1:0] s_574;
  wire [0:0] s_575;
  wire [0:0] s_576;
  wire [0:0] s_577;
  wire [0:0] s_578;
  wire [0:0] s_579;
  wire [0:0] s_580;
  wire [1:0] s_581;
  wire [0:0] s_582;
  wire [0:0] s_583;
  wire [0:0] s_584;
  wire [0:0] s_585;
  wire [0:0] s_586;
  wire [0:0] s_587;
  wire [2:0] s_588;
  wire [0:0] s_589;
  wire [0:0] s_590;
  wire [1:0] s_591;
  wire [0:0] s_592;
  wire [0:0] s_593;
  wire [0:0] s_594;
  wire [1:0] s_595;
  wire [3:0] s_596;
  wire [0:0] s_597;
  wire [0:0] s_598;
  wire [0:0] s_599;
  wire [0:0] s_600;
  wire [0:0] s_601;
  wire [0:0] s_602;
  wire [0:0] s_603;
  wire [1:0] s_604;
  wire [0:0] s_605;
  wire [0:0] s_606;
  wire [0:0] s_607;
  wire [1:0] s_608;
  wire [0:0] s_609;
  wire [0:0] s_610;
  wire [0:0] s_611;
  wire [0:0] s_612;
  wire [0:0] s_613;
  wire [0:0] s_614;
  wire [1:0] s_615;
  wire [0:0] s_616;
  wire [0:0] s_617;
  wire [0:0] s_618;
  wire [0:0] s_619;
  wire [0:0] s_620;
  wire [2:0] s_621;
  wire [0:0] s_622;
  wire [0:0] s_623;
  wire [1:0] s_624;
  wire [1:0] s_625;
  wire [1:0] s_626;
  wire [0:0] s_627;
  wire [3:0] s_628;
  wire [0:0] s_629;
  wire [0:0] s_630;
  wire [2:0] s_631;
  wire [0:0] s_632;
  wire [0:0] s_633;
  wire [1:0] s_634;
  wire [0:0] s_635;
  wire [0:0] s_636;
  wire [0:0] s_637;
  wire [1:0] s_638;
  wire [3:0] s_639;
  wire [7:0] s_640;
  wire [0:0] s_641;
  wire [0:0] s_642;
  wire [0:0] s_643;
  wire [0:0] s_644;
  wire [0:0] s_645;
  wire [0:0] s_646;
  wire [0:0] s_647;
  wire [1:0] s_648;
  wire [0:0] s_649;
  wire [0:0] s_650;
  wire [0:0] s_651;
  wire [1:0] s_652;
  wire [0:0] s_653;
  wire [0:0] s_654;
  wire [0:0] s_655;
  wire [0:0] s_656;
  wire [0:0] s_657;
  wire [0:0] s_658;
  wire [1:0] s_659;
  wire [0:0] s_660;
  wire [0:0] s_661;
  wire [0:0] s_662;
  wire [0:0] s_663;
  wire [0:0] s_664;
  wire [0:0] s_665;
  wire [2:0] s_666;
  wire [0:0] s_667;
  wire [0:0] s_668;
  wire [1:0] s_669;
  wire [0:0] s_670;
  wire [0:0] s_671;
  wire [0:0] s_672;
  wire [1:0] s_673;
  wire [3:0] s_674;
  wire [0:0] s_675;
  wire [0:0] s_676;
  wire [0:0] s_677;
  wire [0:0] s_678;
  wire [0:0] s_679;
  wire [0:0] s_680;
  wire [0:0] s_681;
  wire [1:0] s_682;
  wire [0:0] s_683;
  wire [0:0] s_684;
  wire [0:0] s_685;
  wire [1:0] s_686;
  wire [0:0] s_687;
  wire [0:0] s_688;
  wire [0:0] s_689;
  wire [0:0] s_690;
  wire [0:0] s_691;
  wire [0:0] s_692;
  wire [1:0] s_693;
  wire [0:0] s_694;
  wire [0:0] s_695;
  wire [0:0] s_696;
  wire [0:0] s_697;
  wire [0:0] s_698;
  wire [2:0] s_699;
  wire [0:0] s_700;
  wire [0:0] s_701;
  wire [1:0] s_702;
  wire [1:0] s_703;
  wire [1:0] s_704;
  wire [3:0] s_705;
  wire [0:0] s_706;
  wire [0:0] s_707;
  wire [2:0] s_708;
  wire [2:0] s_709;
  wire [2:0] s_710;
  wire [0:0] s_711;
  wire [4:0] s_712;
  wire [0:0] s_713;
  wire [0:0] s_714;
  wire [3:0] s_715;
  wire [0:0] s_716;
  wire [0:0] s_717;
  wire [2:0] s_718;
  wire [0:0] s_719;
  wire [0:0] s_720;
  wire [1:0] s_721;
  wire [0:0] s_722;
  wire [0:0] s_723;
  wire [0:0] s_724;
  wire [1:0] s_725;
  wire [3:0] s_726;
  wire [7:0] s_727;
  wire [15:0] s_728;
  wire [0:0] s_729;
  wire [0:0] s_730;
  wire [0:0] s_731;
  wire [0:0] s_732;
  wire [0:0] s_733;
  wire [0:0] s_734;
  wire [0:0] s_735;
  wire [1:0] s_736;
  wire [0:0] s_737;
  wire [0:0] s_738;
  wire [0:0] s_739;
  wire [1:0] s_740;
  wire [0:0] s_741;
  wire [0:0] s_742;
  wire [0:0] s_743;
  wire [0:0] s_744;
  wire [0:0] s_745;
  wire [0:0] s_746;
  wire [1:0] s_747;
  wire [0:0] s_748;
  wire [0:0] s_749;
  wire [0:0] s_750;
  wire [0:0] s_751;
  wire [0:0] s_752;
  wire [0:0] s_753;
  wire [2:0] s_754;
  wire [0:0] s_755;
  wire [0:0] s_756;
  wire [1:0] s_757;
  wire [0:0] s_758;
  wire [0:0] s_759;
  wire [0:0] s_760;
  wire [1:0] s_761;
  wire [3:0] s_762;
  wire [0:0] s_763;
  wire [0:0] s_764;
  wire [0:0] s_765;
  wire [0:0] s_766;
  wire [0:0] s_767;
  wire [0:0] s_768;
  wire [0:0] s_769;
  wire [1:0] s_770;
  wire [0:0] s_771;
  wire [0:0] s_772;
  wire [0:0] s_773;
  wire [1:0] s_774;
  wire [0:0] s_775;
  wire [0:0] s_776;
  wire [0:0] s_777;
  wire [0:0] s_778;
  wire [0:0] s_779;
  wire [0:0] s_780;
  wire [1:0] s_781;
  wire [0:0] s_782;
  wire [0:0] s_783;
  wire [0:0] s_784;
  wire [0:0] s_785;
  wire [0:0] s_786;
  wire [2:0] s_787;
  wire [0:0] s_788;
  wire [0:0] s_789;
  wire [1:0] s_790;
  wire [1:0] s_791;
  wire [1:0] s_792;
  wire [0:0] s_793;
  wire [3:0] s_794;
  wire [0:0] s_795;
  wire [0:0] s_796;
  wire [2:0] s_797;
  wire [0:0] s_798;
  wire [0:0] s_799;
  wire [1:0] s_800;
  wire [0:0] s_801;
  wire [0:0] s_802;
  wire [0:0] s_803;
  wire [1:0] s_804;
  wire [3:0] s_805;
  wire [7:0] s_806;
  wire [0:0] s_807;
  wire [0:0] s_808;
  wire [0:0] s_809;
  wire [0:0] s_810;
  wire [0:0] s_811;
  wire [0:0] s_812;
  wire [0:0] s_813;
  wire [1:0] s_814;
  wire [0:0] s_815;
  wire [0:0] s_816;
  wire [0:0] s_817;
  wire [1:0] s_818;
  wire [0:0] s_819;
  wire [0:0] s_820;
  wire [0:0] s_821;
  wire [0:0] s_822;
  wire [0:0] s_823;
  wire [0:0] s_824;
  wire [1:0] s_825;
  wire [0:0] s_826;
  wire [0:0] s_827;
  wire [0:0] s_828;
  wire [0:0] s_829;
  wire [0:0] s_830;
  wire [0:0] s_831;
  wire [2:0] s_832;
  wire [0:0] s_833;
  wire [0:0] s_834;
  wire [1:0] s_835;
  wire [0:0] s_836;
  wire [0:0] s_837;
  wire [0:0] s_838;
  wire [1:0] s_839;
  wire [3:0] s_840;
  wire [0:0] s_841;
  wire [0:0] s_842;
  wire [0:0] s_843;
  wire [0:0] s_844;
  wire [0:0] s_845;
  wire [0:0] s_846;
  wire [0:0] s_847;
  wire [1:0] s_848;
  wire [0:0] s_849;
  wire [0:0] s_850;
  wire [0:0] s_851;
  wire [1:0] s_852;
  wire [0:0] s_853;
  wire [0:0] s_854;
  wire [0:0] s_855;
  wire [0:0] s_856;
  wire [0:0] s_857;
  wire [0:0] s_858;
  wire [1:0] s_859;
  wire [0:0] s_860;
  wire [0:0] s_861;
  wire [0:0] s_862;
  wire [0:0] s_863;
  wire [0:0] s_864;
  wire [2:0] s_865;
  wire [0:0] s_866;
  wire [0:0] s_867;
  wire [1:0] s_868;
  wire [1:0] s_869;
  wire [1:0] s_870;
  wire [3:0] s_871;
  wire [0:0] s_872;
  wire [0:0] s_873;
  wire [2:0] s_874;
  wire [2:0] s_875;
  wire [2:0] s_876;
  wire [4:0] s_877;
  wire [0:0] s_878;
  wire [0:0] s_879;
  wire [3:0] s_880;
  wire [3:0] s_881;
  wire [3:0] s_882;
  wire [5:0] s_883;
  wire [0:0] s_884;
  wire [0:0] s_885;
  wire [4:0] s_886;
  wire [4:0] s_887;
  wire [4:0] s_888;
  wire [12:0] s_889;
  wire [12:0] s_890;
  wire [12:0] s_891;
  wire [10:0] s_892;
  wire [10:0] s_893;
  wire [12:0] s_894;
  wire [0:0] s_895;
  wire [12:0] s_896;
  wire [12:0] s_897;
  wire [0:0] s_898;
  wire [0:0] s_899;
  wire [12:0] s_900;
  wire [12:0] s_901;
  wire [12:0] s_902;
  wire [5:0] s_903;
  wire [108:0] s_904;
  wire [0:0] s_905;
  wire [109:0] s_906;
  wire [109:0] s_907;
  wire [109:0] s_908;
  wire [109:0] s_909;
  wire [108:0] s_910;
  wire [5:0] s_911;
  wire [106:0] s_912;
  wire [108:0] s_913;
  wire [0:0] s_914;
  wire [109:0] s_915;
  wire [109:0] s_916;
  wire [109:0] s_917;
  wire [108:0] s_918;
  wire [5:0] s_919;
  wire [104:0] s_920;
  wire [108:0] s_921;
  wire [0:0] s_922;
  wire [109:0] s_923;
  wire [109:0] s_924;
  wire [109:0] s_925;
  wire [108:0] s_926;
  wire [5:0] s_927;
  wire [102:0] s_928;
  wire [108:0] s_929;
  wire [0:0] s_930;
  wire [109:0] s_931;
  wire [109:0] s_932;
  wire [109:0] s_933;
  wire [108:0] s_934;
  wire [5:0] s_935;
  wire [100:0] s_936;
  wire [108:0] s_937;
  wire [0:0] s_938;
  wire [109:0] s_939;
  wire [109:0] s_940;
  wire [109:0] s_941;
  wire [108:0] s_942;
  wire [5:0] s_943;
  wire [98:0] s_944;
  wire [108:0] s_945;
  wire [0:0] s_946;
  wire [109:0] s_947;
  wire [109:0] s_948;
  wire [109:0] s_949;
  wire [108:0] s_950;
  wire [5:0] s_951;
  wire [96:0] s_952;
  wire [108:0] s_953;
  wire [0:0] s_954;
  wire [109:0] s_955;
  wire [109:0] s_956;
  wire [109:0] s_957;
  wire [108:0] s_958;
  wire [5:0] s_959;
  wire [94:0] s_960;
  wire [108:0] s_961;
  wire [0:0] s_962;
  wire [109:0] s_963;
  wire [109:0] s_964;
  wire [109:0] s_965;
  wire [108:0] s_966;
  wire [5:0] s_967;
  wire [92:0] s_968;
  wire [108:0] s_969;
  wire [0:0] s_970;
  wire [109:0] s_971;
  wire [109:0] s_972;
  wire [109:0] s_973;
  wire [108:0] s_974;
  wire [5:0] s_975;
  wire [90:0] s_976;
  wire [108:0] s_977;
  wire [0:0] s_978;
  wire [109:0] s_979;
  wire [109:0] s_980;
  wire [109:0] s_981;
  wire [108:0] s_982;
  wire [5:0] s_983;
  wire [88:0] s_984;
  wire [108:0] s_985;
  wire [0:0] s_986;
  wire [109:0] s_987;
  wire [109:0] s_988;
  wire [109:0] s_989;
  wire [108:0] s_990;
  wire [5:0] s_991;
  wire [86:0] s_992;
  wire [108:0] s_993;
  wire [0:0] s_994;
  wire [109:0] s_995;
  wire [109:0] s_996;
  wire [109:0] s_997;
  wire [108:0] s_998;
  wire [5:0] s_999;
  wire [84:0] s_1000;
  wire [108:0] s_1001;
  wire [0:0] s_1002;
  wire [109:0] s_1003;
  wire [109:0] s_1004;
  wire [109:0] s_1005;
  wire [108:0] s_1006;
  wire [5:0] s_1007;
  wire [82:0] s_1008;
  wire [108:0] s_1009;
  wire [0:0] s_1010;
  wire [109:0] s_1011;
  wire [109:0] s_1012;
  wire [109:0] s_1013;
  wire [108:0] s_1014;
  wire [5:0] s_1015;
  wire [80:0] s_1016;
  wire [108:0] s_1017;
  wire [0:0] s_1018;
  wire [109:0] s_1019;
  wire [109:0] s_1020;
  wire [109:0] s_1021;
  wire [108:0] s_1022;
  wire [5:0] s_1023;
  wire [78:0] s_1024;
  wire [108:0] s_1025;
  wire [0:0] s_1026;
  wire [109:0] s_1027;
  wire [109:0] s_1028;
  wire [109:0] s_1029;
  wire [108:0] s_1030;
  wire [5:0] s_1031;
  wire [76:0] s_1032;
  wire [108:0] s_1033;
  wire [0:0] s_1034;
  wire [109:0] s_1035;
  wire [109:0] s_1036;
  wire [109:0] s_1037;
  wire [108:0] s_1038;
  wire [5:0] s_1039;
  wire [74:0] s_1040;
  wire [108:0] s_1041;
  wire [0:0] s_1042;
  wire [109:0] s_1043;
  wire [109:0] s_1044;
  wire [109:0] s_1045;
  wire [108:0] s_1046;
  wire [5:0] s_1047;
  wire [72:0] s_1048;
  wire [108:0] s_1049;
  wire [0:0] s_1050;
  wire [109:0] s_1051;
  wire [109:0] s_1052;
  wire [109:0] s_1053;
  wire [108:0] s_1054;
  wire [5:0] s_1055;
  wire [70:0] s_1056;
  wire [108:0] s_1057;
  wire [0:0] s_1058;
  wire [109:0] s_1059;
  wire [109:0] s_1060;
  wire [109:0] s_1061;
  wire [108:0] s_1062;
  wire [5:0] s_1063;
  wire [68:0] s_1064;
  wire [108:0] s_1065;
  wire [0:0] s_1066;
  wire [109:0] s_1067;
  wire [109:0] s_1068;
  wire [109:0] s_1069;
  wire [108:0] s_1070;
  wire [5:0] s_1071;
  wire [66:0] s_1072;
  wire [108:0] s_1073;
  wire [0:0] s_1074;
  wire [109:0] s_1075;
  wire [109:0] s_1076;
  wire [109:0] s_1077;
  wire [108:0] s_1078;
  wire [5:0] s_1079;
  wire [64:0] s_1080;
  wire [108:0] s_1081;
  wire [0:0] s_1082;
  wire [109:0] s_1083;
  wire [109:0] s_1084;
  wire [109:0] s_1085;
  wire [108:0] s_1086;
  wire [5:0] s_1087;
  wire [62:0] s_1088;
  wire [108:0] s_1089;
  wire [0:0] s_1090;
  wire [109:0] s_1091;
  wire [109:0] s_1092;
  wire [109:0] s_1093;
  wire [108:0] s_1094;
  wire [4:0] s_1095;
  wire [60:0] s_1096;
  wire [108:0] s_1097;
  wire [0:0] s_1098;
  wire [109:0] s_1099;
  wire [109:0] s_1100;
  wire [109:0] s_1101;
  wire [108:0] s_1102;
  wire [4:0] s_1103;
  wire [58:0] s_1104;
  wire [108:0] s_1105;
  wire [0:0] s_1106;
  wire [109:0] s_1107;
  wire [109:0] s_1108;
  wire [109:0] s_1109;
  wire [108:0] s_1110;
  wire [4:0] s_1111;
  wire [56:0] s_1112;
  wire [108:0] s_1113;
  wire [0:0] s_1114;
  wire [109:0] s_1115;
  wire [109:0] s_1116;
  wire [109:0] s_1117;
  wire [108:0] s_1118;
  wire [4:0] s_1119;
  wire [54:0] s_1120;
  wire [108:0] s_1121;
  wire [0:0] s_1122;
  wire [109:0] s_1123;
  wire [109:0] s_1124;
  wire [109:0] s_1125;
  wire [108:0] s_1126;
  wire [4:0] s_1127;
  wire [52:0] s_1128;
  wire [108:0] s_1129;
  wire [0:0] s_1130;
  wire [109:0] s_1131;
  wire [109:0] s_1132;
  wire [109:0] s_1133;
  wire [108:0] s_1134;
  wire [4:0] s_1135;
  wire [50:0] s_1136;
  wire [108:0] s_1137;
  wire [0:0] s_1138;
  wire [109:0] s_1139;
  wire [109:0] s_1140;
  wire [109:0] s_1141;
  wire [108:0] s_1142;
  wire [4:0] s_1143;
  wire [48:0] s_1144;
  wire [108:0] s_1145;
  wire [0:0] s_1146;
  wire [109:0] s_1147;
  wire [109:0] s_1148;
  wire [109:0] s_1149;
  wire [108:0] s_1150;
  wire [4:0] s_1151;
  wire [46:0] s_1152;
  wire [108:0] s_1153;
  wire [0:0] s_1154;
  wire [109:0] s_1155;
  wire [109:0] s_1156;
  wire [109:0] s_1157;
  wire [108:0] s_1158;
  wire [4:0] s_1159;
  wire [44:0] s_1160;
  wire [108:0] s_1161;
  wire [0:0] s_1162;
  wire [109:0] s_1163;
  wire [109:0] s_1164;
  wire [109:0] s_1165;
  wire [108:0] s_1166;
  wire [4:0] s_1167;
  wire [42:0] s_1168;
  wire [108:0] s_1169;
  wire [0:0] s_1170;
  wire [109:0] s_1171;
  wire [109:0] s_1172;
  wire [109:0] s_1173;
  wire [108:0] s_1174;
  wire [4:0] s_1175;
  wire [40:0] s_1176;
  wire [108:0] s_1177;
  wire [0:0] s_1178;
  wire [109:0] s_1179;
  wire [109:0] s_1180;
  wire [109:0] s_1181;
  wire [108:0] s_1182;
  wire [4:0] s_1183;
  wire [38:0] s_1184;
  wire [108:0] s_1185;
  wire [0:0] s_1186;
  wire [109:0] s_1187;
  wire [109:0] s_1188;
  wire [109:0] s_1189;
  wire [108:0] s_1190;
  wire [4:0] s_1191;
  wire [36:0] s_1192;
  wire [108:0] s_1193;
  wire [0:0] s_1194;
  wire [109:0] s_1195;
  wire [109:0] s_1196;
  wire [109:0] s_1197;
  wire [108:0] s_1198;
  wire [4:0] s_1199;
  wire [34:0] s_1200;
  wire [108:0] s_1201;
  wire [0:0] s_1202;
  wire [109:0] s_1203;
  wire [109:0] s_1204;
  wire [109:0] s_1205;
  wire [108:0] s_1206;
  wire [4:0] s_1207;
  wire [32:0] s_1208;
  wire [108:0] s_1209;
  wire [0:0] s_1210;
  wire [109:0] s_1211;
  wire [109:0] s_1212;
  wire [109:0] s_1213;
  wire [108:0] s_1214;
  wire [4:0] s_1215;
  wire [30:0] s_1216;
  wire [108:0] s_1217;
  wire [0:0] s_1218;
  wire [109:0] s_1219;
  wire [109:0] s_1220;
  wire [109:0] s_1221;
  wire [108:0] s_1222;
  wire [3:0] s_1223;
  wire [28:0] s_1224;
  wire [108:0] s_1225;
  wire [0:0] s_1226;
  wire [109:0] s_1227;
  wire [109:0] s_1228;
  wire [109:0] s_1229;
  wire [108:0] s_1230;
  wire [3:0] s_1231;
  wire [26:0] s_1232;
  wire [108:0] s_1233;
  wire [0:0] s_1234;
  wire [109:0] s_1235;
  wire [109:0] s_1236;
  wire [109:0] s_1237;
  wire [108:0] s_1238;
  wire [3:0] s_1239;
  wire [24:0] s_1240;
  wire [108:0] s_1241;
  wire [0:0] s_1242;
  wire [109:0] s_1243;
  wire [109:0] s_1244;
  wire [109:0] s_1245;
  wire [108:0] s_1246;
  wire [3:0] s_1247;
  wire [22:0] s_1248;
  wire [108:0] s_1249;
  wire [0:0] s_1250;
  wire [109:0] s_1251;
  wire [109:0] s_1252;
  wire [109:0] s_1253;
  wire [108:0] s_1254;
  wire [3:0] s_1255;
  wire [20:0] s_1256;
  wire [108:0] s_1257;
  wire [0:0] s_1258;
  wire [109:0] s_1259;
  wire [109:0] s_1260;
  wire [109:0] s_1261;
  wire [108:0] s_1262;
  wire [3:0] s_1263;
  wire [18:0] s_1264;
  wire [108:0] s_1265;
  wire [0:0] s_1266;
  wire [109:0] s_1267;
  wire [109:0] s_1268;
  wire [109:0] s_1269;
  wire [108:0] s_1270;
  wire [3:0] s_1271;
  wire [16:0] s_1272;
  wire [108:0] s_1273;
  wire [0:0] s_1274;
  wire [109:0] s_1275;
  wire [109:0] s_1276;
  wire [109:0] s_1277;
  wire [108:0] s_1278;
  wire [3:0] s_1279;
  wire [14:0] s_1280;
  wire [108:0] s_1281;
  wire [0:0] s_1282;
  wire [109:0] s_1283;
  wire [109:0] s_1284;
  wire [109:0] s_1285;
  wire [108:0] s_1286;
  wire [2:0] s_1287;
  wire [12:0] s_1288;
  wire [108:0] s_1289;
  wire [0:0] s_1290;
  wire [109:0] s_1291;
  wire [109:0] s_1292;
  wire [109:0] s_1293;
  wire [108:0] s_1294;
  wire [2:0] s_1295;
  wire [10:0] s_1296;
  wire [108:0] s_1297;
  wire [0:0] s_1298;
  wire [109:0] s_1299;
  wire [109:0] s_1300;
  wire [109:0] s_1301;
  wire [108:0] s_1302;
  wire [2:0] s_1303;
  wire [8:0] s_1304;
  wire [108:0] s_1305;
  wire [0:0] s_1306;
  wire [109:0] s_1307;
  wire [109:0] s_1308;
  wire [109:0] s_1309;
  wire [108:0] s_1310;
  wire [2:0] s_1311;
  wire [6:0] s_1312;
  wire [108:0] s_1313;
  wire [0:0] s_1314;
  wire [109:0] s_1315;
  wire [109:0] s_1316;
  wire [109:0] s_1317;
  wire [108:0] s_1318;
  wire [1:0] s_1319;
  wire [4:0] s_1320;
  wire [108:0] s_1321;
  wire [0:0] s_1322;
  wire [109:0] s_1323;
  wire [109:0] s_1324;
  wire [109:0] s_1325;
  wire [108:0] s_1326;
  wire [1:0] s_1327;
  wire [2:0] s_1328;
  wire [108:0] s_1329;
  wire [0:0] s_1330;
  wire [109:0] s_1331;
  wire [109:0] s_1332;
  wire [109:0] s_1333;
  wire [108:0] s_1334;
  wire [0:0] s_1335;
  wire [0:0] s_1336;
  wire [12:0] s_1337;
  wire [12:0] s_1338;
  wire [0:0] s_1339;
  wire [12:0] s_1340;
  wire [12:0] s_1341;
  wire [12:0] s_1342;
  wire [12:0] s_1343;
  wire [12:0] s_1344;
  wire [12:0] s_1345;
  wire [0:0] s_1346;
  wire [12:0] s_1347;
  wire [0:0] s_1348;
  wire [12:0] s_1349;
  wire [12:0] s_1350;
  wire [6:0] s_1351;
  wire [6:0] s_1352;
  wire [0:0] s_1353;
  wire [0:0] s_1354;
  wire [5:0] s_1355;
  wire [0:0] s_1356;
  wire [0:0] s_1357;
  wire [4:0] s_1358;
  wire [0:0] s_1359;
  wire [0:0] s_1360;
  wire [3:0] s_1361;
  wire [0:0] s_1362;
  wire [0:0] s_1363;
  wire [2:0] s_1364;
  wire [0:0] s_1365;
  wire [0:0] s_1366;
  wire [1:0] s_1367;
  wire [0:0] s_1368;
  wire [0:0] s_1369;
  wire [0:0] s_1370;
  wire [1:0] s_1371;
  wire [3:0] s_1372;
  wire [7:0] s_1373;
  wire [15:0] s_1374;
  wire [31:0] s_1375;
  wire [63:0] s_1376;
  wire [62:0] s_1377;
  wire [61:0] s_1378;
  wire [60:0] s_1379;
  wire [59:0] s_1380;
  wire [58:0] s_1381;
  wire [57:0] s_1382;
  wire [56:0] s_1383;
  wire [55:0] s_1384;
  wire [54:0] s_1385;
  wire [0:0] s_1386;
  wire [0:0] s_1387;
  wire [0:0] s_1388;
  wire [0:0] s_1389;
  wire [0:0] s_1390;
  wire [0:0] s_1391;
  wire [0:0] s_1392;
  wire [0:0] s_1393;
  wire [0:0] s_1394;
  wire [0:0] s_1395;
  wire [0:0] s_1396;
  wire [0:0] s_1397;
  wire [0:0] s_1398;
  wire [0:0] s_1399;
  wire [0:0] s_1400;
  wire [0:0] s_1401;
  wire [0:0] s_1402;
  wire [1:0] s_1403;
  wire [0:0] s_1404;
  wire [0:0] s_1405;
  wire [0:0] s_1406;
  wire [1:0] s_1407;
  wire [0:0] s_1408;
  wire [0:0] s_1409;
  wire [0:0] s_1410;
  wire [0:0] s_1411;
  wire [0:0] s_1412;
  wire [0:0] s_1413;
  wire [1:0] s_1414;
  wire [0:0] s_1415;
  wire [0:0] s_1416;
  wire [0:0] s_1417;
  wire [0:0] s_1418;
  wire [0:0] s_1419;
  wire [0:0] s_1420;
  wire [2:0] s_1421;
  wire [0:0] s_1422;
  wire [0:0] s_1423;
  wire [1:0] s_1424;
  wire [0:0] s_1425;
  wire [0:0] s_1426;
  wire [0:0] s_1427;
  wire [1:0] s_1428;
  wire [3:0] s_1429;
  wire [0:0] s_1430;
  wire [0:0] s_1431;
  wire [0:0] s_1432;
  wire [0:0] s_1433;
  wire [0:0] s_1434;
  wire [0:0] s_1435;
  wire [0:0] s_1436;
  wire [1:0] s_1437;
  wire [0:0] s_1438;
  wire [0:0] s_1439;
  wire [0:0] s_1440;
  wire [1:0] s_1441;
  wire [0:0] s_1442;
  wire [0:0] s_1443;
  wire [0:0] s_1444;
  wire [0:0] s_1445;
  wire [0:0] s_1446;
  wire [0:0] s_1447;
  wire [1:0] s_1448;
  wire [0:0] s_1449;
  wire [0:0] s_1450;
  wire [0:0] s_1451;
  wire [0:0] s_1452;
  wire [0:0] s_1453;
  wire [2:0] s_1454;
  wire [0:0] s_1455;
  wire [0:0] s_1456;
  wire [1:0] s_1457;
  wire [1:0] s_1458;
  wire [1:0] s_1459;
  wire [0:0] s_1460;
  wire [3:0] s_1461;
  wire [0:0] s_1462;
  wire [0:0] s_1463;
  wire [2:0] s_1464;
  wire [0:0] s_1465;
  wire [0:0] s_1466;
  wire [1:0] s_1467;
  wire [0:0] s_1468;
  wire [0:0] s_1469;
  wire [0:0] s_1470;
  wire [1:0] s_1471;
  wire [3:0] s_1472;
  wire [7:0] s_1473;
  wire [0:0] s_1474;
  wire [0:0] s_1475;
  wire [0:0] s_1476;
  wire [0:0] s_1477;
  wire [0:0] s_1478;
  wire [0:0] s_1479;
  wire [0:0] s_1480;
  wire [1:0] s_1481;
  wire [0:0] s_1482;
  wire [0:0] s_1483;
  wire [0:0] s_1484;
  wire [1:0] s_1485;
  wire [0:0] s_1486;
  wire [0:0] s_1487;
  wire [0:0] s_1488;
  wire [0:0] s_1489;
  wire [0:0] s_1490;
  wire [0:0] s_1491;
  wire [1:0] s_1492;
  wire [0:0] s_1493;
  wire [0:0] s_1494;
  wire [0:0] s_1495;
  wire [0:0] s_1496;
  wire [0:0] s_1497;
  wire [0:0] s_1498;
  wire [2:0] s_1499;
  wire [0:0] s_1500;
  wire [0:0] s_1501;
  wire [1:0] s_1502;
  wire [0:0] s_1503;
  wire [0:0] s_1504;
  wire [0:0] s_1505;
  wire [1:0] s_1506;
  wire [3:0] s_1507;
  wire [0:0] s_1508;
  wire [0:0] s_1509;
  wire [0:0] s_1510;
  wire [0:0] s_1511;
  wire [0:0] s_1512;
  wire [0:0] s_1513;
  wire [0:0] s_1514;
  wire [1:0] s_1515;
  wire [0:0] s_1516;
  wire [0:0] s_1517;
  wire [0:0] s_1518;
  wire [1:0] s_1519;
  wire [0:0] s_1520;
  wire [0:0] s_1521;
  wire [0:0] s_1522;
  wire [0:0] s_1523;
  wire [0:0] s_1524;
  wire [0:0] s_1525;
  wire [1:0] s_1526;
  wire [0:0] s_1527;
  wire [0:0] s_1528;
  wire [0:0] s_1529;
  wire [0:0] s_1530;
  wire [0:0] s_1531;
  wire [2:0] s_1532;
  wire [0:0] s_1533;
  wire [0:0] s_1534;
  wire [1:0] s_1535;
  wire [1:0] s_1536;
  wire [1:0] s_1537;
  wire [3:0] s_1538;
  wire [0:0] s_1539;
  wire [0:0] s_1540;
  wire [2:0] s_1541;
  wire [2:0] s_1542;
  wire [2:0] s_1543;
  wire [0:0] s_1544;
  wire [4:0] s_1545;
  wire [0:0] s_1546;
  wire [0:0] s_1547;
  wire [3:0] s_1548;
  wire [0:0] s_1549;
  wire [0:0] s_1550;
  wire [2:0] s_1551;
  wire [0:0] s_1552;
  wire [0:0] s_1553;
  wire [1:0] s_1554;
  wire [0:0] s_1555;
  wire [0:0] s_1556;
  wire [0:0] s_1557;
  wire [1:0] s_1558;
  wire [3:0] s_1559;
  wire [7:0] s_1560;
  wire [15:0] s_1561;
  wire [0:0] s_1562;
  wire [0:0] s_1563;
  wire [0:0] s_1564;
  wire [0:0] s_1565;
  wire [0:0] s_1566;
  wire [0:0] s_1567;
  wire [0:0] s_1568;
  wire [1:0] s_1569;
  wire [0:0] s_1570;
  wire [0:0] s_1571;
  wire [0:0] s_1572;
  wire [1:0] s_1573;
  wire [0:0] s_1574;
  wire [0:0] s_1575;
  wire [0:0] s_1576;
  wire [0:0] s_1577;
  wire [0:0] s_1578;
  wire [0:0] s_1579;
  wire [1:0] s_1580;
  wire [0:0] s_1581;
  wire [0:0] s_1582;
  wire [0:0] s_1583;
  wire [0:0] s_1584;
  wire [0:0] s_1585;
  wire [0:0] s_1586;
  wire [2:0] s_1587;
  wire [0:0] s_1588;
  wire [0:0] s_1589;
  wire [1:0] s_1590;
  wire [0:0] s_1591;
  wire [0:0] s_1592;
  wire [0:0] s_1593;
  wire [1:0] s_1594;
  wire [3:0] s_1595;
  wire [0:0] s_1596;
  wire [0:0] s_1597;
  wire [0:0] s_1598;
  wire [0:0] s_1599;
  wire [0:0] s_1600;
  wire [0:0] s_1601;
  wire [0:0] s_1602;
  wire [1:0] s_1603;
  wire [0:0] s_1604;
  wire [0:0] s_1605;
  wire [0:0] s_1606;
  wire [1:0] s_1607;
  wire [0:0] s_1608;
  wire [0:0] s_1609;
  wire [0:0] s_1610;
  wire [0:0] s_1611;
  wire [0:0] s_1612;
  wire [0:0] s_1613;
  wire [1:0] s_1614;
  wire [0:0] s_1615;
  wire [0:0] s_1616;
  wire [0:0] s_1617;
  wire [0:0] s_1618;
  wire [0:0] s_1619;
  wire [2:0] s_1620;
  wire [0:0] s_1621;
  wire [0:0] s_1622;
  wire [1:0] s_1623;
  wire [1:0] s_1624;
  wire [1:0] s_1625;
  wire [0:0] s_1626;
  wire [3:0] s_1627;
  wire [0:0] s_1628;
  wire [0:0] s_1629;
  wire [2:0] s_1630;
  wire [0:0] s_1631;
  wire [0:0] s_1632;
  wire [1:0] s_1633;
  wire [0:0] s_1634;
  wire [0:0] s_1635;
  wire [0:0] s_1636;
  wire [1:0] s_1637;
  wire [3:0] s_1638;
  wire [7:0] s_1639;
  wire [0:0] s_1640;
  wire [0:0] s_1641;
  wire [0:0] s_1642;
  wire [0:0] s_1643;
  wire [0:0] s_1644;
  wire [0:0] s_1645;
  wire [0:0] s_1646;
  wire [1:0] s_1647;
  wire [0:0] s_1648;
  wire [0:0] s_1649;
  wire [0:0] s_1650;
  wire [1:0] s_1651;
  wire [0:0] s_1652;
  wire [0:0] s_1653;
  wire [0:0] s_1654;
  wire [0:0] s_1655;
  wire [0:0] s_1656;
  wire [0:0] s_1657;
  wire [1:0] s_1658;
  wire [0:0] s_1659;
  wire [0:0] s_1660;
  wire [0:0] s_1661;
  wire [0:0] s_1662;
  wire [0:0] s_1663;
  wire [0:0] s_1664;
  wire [2:0] s_1665;
  wire [0:0] s_1666;
  wire [0:0] s_1667;
  wire [1:0] s_1668;
  wire [0:0] s_1669;
  wire [0:0] s_1670;
  wire [0:0] s_1671;
  wire [1:0] s_1672;
  wire [3:0] s_1673;
  wire [0:0] s_1674;
  wire [0:0] s_1675;
  wire [0:0] s_1676;
  wire [0:0] s_1677;
  wire [0:0] s_1678;
  wire [0:0] s_1679;
  wire [0:0] s_1680;
  wire [1:0] s_1681;
  wire [0:0] s_1682;
  wire [0:0] s_1683;
  wire [0:0] s_1684;
  wire [1:0] s_1685;
  wire [0:0] s_1686;
  wire [0:0] s_1687;
  wire [0:0] s_1688;
  wire [0:0] s_1689;
  wire [0:0] s_1690;
  wire [0:0] s_1691;
  wire [1:0] s_1692;
  wire [0:0] s_1693;
  wire [0:0] s_1694;
  wire [0:0] s_1695;
  wire [0:0] s_1696;
  wire [0:0] s_1697;
  wire [2:0] s_1698;
  wire [0:0] s_1699;
  wire [0:0] s_1700;
  wire [1:0] s_1701;
  wire [1:0] s_1702;
  wire [1:0] s_1703;
  wire [3:0] s_1704;
  wire [0:0] s_1705;
  wire [0:0] s_1706;
  wire [2:0] s_1707;
  wire [2:0] s_1708;
  wire [2:0] s_1709;
  wire [4:0] s_1710;
  wire [0:0] s_1711;
  wire [0:0] s_1712;
  wire [3:0] s_1713;
  wire [3:0] s_1714;
  wire [3:0] s_1715;
  wire [0:0] s_1716;
  wire [5:0] s_1717;
  wire [0:0] s_1718;
  wire [0:0] s_1719;
  wire [4:0] s_1720;
  wire [0:0] s_1721;
  wire [0:0] s_1722;
  wire [3:0] s_1723;
  wire [0:0] s_1724;
  wire [0:0] s_1725;
  wire [2:0] s_1726;
  wire [0:0] s_1727;
  wire [0:0] s_1728;
  wire [1:0] s_1729;
  wire [0:0] s_1730;
  wire [0:0] s_1731;
  wire [0:0] s_1732;
  wire [1:0] s_1733;
  wire [3:0] s_1734;
  wire [7:0] s_1735;
  wire [15:0] s_1736;
  wire [31:0] s_1737;
  wire [0:0] s_1738;
  wire [0:0] s_1739;
  wire [0:0] s_1740;
  wire [0:0] s_1741;
  wire [0:0] s_1742;
  wire [0:0] s_1743;
  wire [0:0] s_1744;
  wire [1:0] s_1745;
  wire [0:0] s_1746;
  wire [0:0] s_1747;
  wire [0:0] s_1748;
  wire [1:0] s_1749;
  wire [0:0] s_1750;
  wire [0:0] s_1751;
  wire [0:0] s_1752;
  wire [0:0] s_1753;
  wire [0:0] s_1754;
  wire [0:0] s_1755;
  wire [1:0] s_1756;
  wire [0:0] s_1757;
  wire [0:0] s_1758;
  wire [0:0] s_1759;
  wire [0:0] s_1760;
  wire [0:0] s_1761;
  wire [0:0] s_1762;
  wire [2:0] s_1763;
  wire [0:0] s_1764;
  wire [0:0] s_1765;
  wire [1:0] s_1766;
  wire [0:0] s_1767;
  wire [0:0] s_1768;
  wire [0:0] s_1769;
  wire [1:0] s_1770;
  wire [3:0] s_1771;
  wire [0:0] s_1772;
  wire [0:0] s_1773;
  wire [0:0] s_1774;
  wire [0:0] s_1775;
  wire [0:0] s_1776;
  wire [0:0] s_1777;
  wire [0:0] s_1778;
  wire [1:0] s_1779;
  wire [0:0] s_1780;
  wire [0:0] s_1781;
  wire [0:0] s_1782;
  wire [1:0] s_1783;
  wire [0:0] s_1784;
  wire [0:0] s_1785;
  wire [0:0] s_1786;
  wire [0:0] s_1787;
  wire [0:0] s_1788;
  wire [0:0] s_1789;
  wire [1:0] s_1790;
  wire [0:0] s_1791;
  wire [0:0] s_1792;
  wire [0:0] s_1793;
  wire [0:0] s_1794;
  wire [0:0] s_1795;
  wire [2:0] s_1796;
  wire [0:0] s_1797;
  wire [0:0] s_1798;
  wire [1:0] s_1799;
  wire [1:0] s_1800;
  wire [1:0] s_1801;
  wire [0:0] s_1802;
  wire [3:0] s_1803;
  wire [0:0] s_1804;
  wire [0:0] s_1805;
  wire [2:0] s_1806;
  wire [0:0] s_1807;
  wire [0:0] s_1808;
  wire [1:0] s_1809;
  wire [0:0] s_1810;
  wire [0:0] s_1811;
  wire [0:0] s_1812;
  wire [1:0] s_1813;
  wire [3:0] s_1814;
  wire [7:0] s_1815;
  wire [0:0] s_1816;
  wire [0:0] s_1817;
  wire [0:0] s_1818;
  wire [0:0] s_1819;
  wire [0:0] s_1820;
  wire [0:0] s_1821;
  wire [0:0] s_1822;
  wire [1:0] s_1823;
  wire [0:0] s_1824;
  wire [0:0] s_1825;
  wire [0:0] s_1826;
  wire [1:0] s_1827;
  wire [0:0] s_1828;
  wire [0:0] s_1829;
  wire [0:0] s_1830;
  wire [0:0] s_1831;
  wire [0:0] s_1832;
  wire [0:0] s_1833;
  wire [1:0] s_1834;
  wire [0:0] s_1835;
  wire [0:0] s_1836;
  wire [0:0] s_1837;
  wire [0:0] s_1838;
  wire [0:0] s_1839;
  wire [0:0] s_1840;
  wire [2:0] s_1841;
  wire [0:0] s_1842;
  wire [0:0] s_1843;
  wire [1:0] s_1844;
  wire [0:0] s_1845;
  wire [0:0] s_1846;
  wire [0:0] s_1847;
  wire [1:0] s_1848;
  wire [3:0] s_1849;
  wire [0:0] s_1850;
  wire [0:0] s_1851;
  wire [0:0] s_1852;
  wire [0:0] s_1853;
  wire [0:0] s_1854;
  wire [0:0] s_1855;
  wire [0:0] s_1856;
  wire [1:0] s_1857;
  wire [0:0] s_1858;
  wire [0:0] s_1859;
  wire [0:0] s_1860;
  wire [1:0] s_1861;
  wire [0:0] s_1862;
  wire [0:0] s_1863;
  wire [0:0] s_1864;
  wire [0:0] s_1865;
  wire [0:0] s_1866;
  wire [0:0] s_1867;
  wire [1:0] s_1868;
  wire [0:0] s_1869;
  wire [0:0] s_1870;
  wire [0:0] s_1871;
  wire [0:0] s_1872;
  wire [0:0] s_1873;
  wire [2:0] s_1874;
  wire [0:0] s_1875;
  wire [0:0] s_1876;
  wire [1:0] s_1877;
  wire [1:0] s_1878;
  wire [1:0] s_1879;
  wire [3:0] s_1880;
  wire [0:0] s_1881;
  wire [0:0] s_1882;
  wire [2:0] s_1883;
  wire [2:0] s_1884;
  wire [2:0] s_1885;
  wire [0:0] s_1886;
  wire [4:0] s_1887;
  wire [0:0] s_1888;
  wire [0:0] s_1889;
  wire [3:0] s_1890;
  wire [0:0] s_1891;
  wire [0:0] s_1892;
  wire [2:0] s_1893;
  wire [0:0] s_1894;
  wire [0:0] s_1895;
  wire [1:0] s_1896;
  wire [0:0] s_1897;
  wire [0:0] s_1898;
  wire [0:0] s_1899;
  wire [1:0] s_1900;
  wire [3:0] s_1901;
  wire [7:0] s_1902;
  wire [15:0] s_1903;
  wire [0:0] s_1904;
  wire [0:0] s_1905;
  wire [0:0] s_1906;
  wire [0:0] s_1907;
  wire [0:0] s_1908;
  wire [0:0] s_1909;
  wire [0:0] s_1910;
  wire [1:0] s_1911;
  wire [0:0] s_1912;
  wire [0:0] s_1913;
  wire [0:0] s_1914;
  wire [1:0] s_1915;
  wire [0:0] s_1916;
  wire [0:0] s_1917;
  wire [0:0] s_1918;
  wire [0:0] s_1919;
  wire [0:0] s_1920;
  wire [0:0] s_1921;
  wire [1:0] s_1922;
  wire [0:0] s_1923;
  wire [0:0] s_1924;
  wire [0:0] s_1925;
  wire [0:0] s_1926;
  wire [0:0] s_1927;
  wire [0:0] s_1928;
  wire [2:0] s_1929;
  wire [0:0] s_1930;
  wire [0:0] s_1931;
  wire [1:0] s_1932;
  wire [0:0] s_1933;
  wire [0:0] s_1934;
  wire [0:0] s_1935;
  wire [1:0] s_1936;
  wire [3:0] s_1937;
  wire [0:0] s_1938;
  wire [0:0] s_1939;
  wire [0:0] s_1940;
  wire [0:0] s_1941;
  wire [0:0] s_1942;
  wire [0:0] s_1943;
  wire [0:0] s_1944;
  wire [1:0] s_1945;
  wire [0:0] s_1946;
  wire [0:0] s_1947;
  wire [0:0] s_1948;
  wire [1:0] s_1949;
  wire [0:0] s_1950;
  wire [0:0] s_1951;
  wire [0:0] s_1952;
  wire [0:0] s_1953;
  wire [0:0] s_1954;
  wire [0:0] s_1955;
  wire [1:0] s_1956;
  wire [0:0] s_1957;
  wire [0:0] s_1958;
  wire [0:0] s_1959;
  wire [0:0] s_1960;
  wire [0:0] s_1961;
  wire [2:0] s_1962;
  wire [0:0] s_1963;
  wire [0:0] s_1964;
  wire [1:0] s_1965;
  wire [1:0] s_1966;
  wire [1:0] s_1967;
  wire [0:0] s_1968;
  wire [3:0] s_1969;
  wire [0:0] s_1970;
  wire [0:0] s_1971;
  wire [2:0] s_1972;
  wire [0:0] s_1973;
  wire [0:0] s_1974;
  wire [1:0] s_1975;
  wire [0:0] s_1976;
  wire [0:0] s_1977;
  wire [0:0] s_1978;
  wire [1:0] s_1979;
  wire [3:0] s_1980;
  wire [7:0] s_1981;
  wire [0:0] s_1982;
  wire [0:0] s_1983;
  wire [0:0] s_1984;
  wire [0:0] s_1985;
  wire [0:0] s_1986;
  wire [0:0] s_1987;
  wire [0:0] s_1988;
  wire [1:0] s_1989;
  wire [0:0] s_1990;
  wire [0:0] s_1991;
  wire [0:0] s_1992;
  wire [1:0] s_1993;
  wire [0:0] s_1994;
  wire [0:0] s_1995;
  wire [0:0] s_1996;
  wire [0:0] s_1997;
  wire [0:0] s_1998;
  wire [0:0] s_1999;
  wire [1:0] s_2000;
  wire [0:0] s_2001;
  wire [0:0] s_2002;
  wire [0:0] s_2003;
  wire [0:0] s_2004;
  wire [0:0] s_2005;
  wire [0:0] s_2006;
  wire [2:0] s_2007;
  wire [0:0] s_2008;
  wire [0:0] s_2009;
  wire [1:0] s_2010;
  wire [0:0] s_2011;
  wire [0:0] s_2012;
  wire [0:0] s_2013;
  wire [1:0] s_2014;
  wire [3:0] s_2015;
  wire [0:0] s_2016;
  wire [0:0] s_2017;
  wire [0:0] s_2018;
  wire [0:0] s_2019;
  wire [0:0] s_2020;
  wire [0:0] s_2021;
  wire [0:0] s_2022;
  wire [1:0] s_2023;
  wire [0:0] s_2024;
  wire [0:0] s_2025;
  wire [0:0] s_2026;
  wire [1:0] s_2027;
  wire [0:0] s_2028;
  wire [0:0] s_2029;
  wire [0:0] s_2030;
  wire [0:0] s_2031;
  wire [0:0] s_2032;
  wire [0:0] s_2033;
  wire [1:0] s_2034;
  wire [0:0] s_2035;
  wire [0:0] s_2036;
  wire [0:0] s_2037;
  wire [0:0] s_2038;
  wire [0:0] s_2039;
  wire [2:0] s_2040;
  wire [0:0] s_2041;
  wire [0:0] s_2042;
  wire [1:0] s_2043;
  wire [1:0] s_2044;
  wire [1:0] s_2045;
  wire [3:0] s_2046;
  wire [0:0] s_2047;
  wire [0:0] s_2048;
  wire [2:0] s_2049;
  wire [2:0] s_2050;
  wire [2:0] s_2051;
  wire [4:0] s_2052;
  wire [0:0] s_2053;
  wire [0:0] s_2054;
  wire [3:0] s_2055;
  wire [3:0] s_2056;
  wire [3:0] s_2057;
  wire [5:0] s_2058;
  wire [0:0] s_2059;
  wire [0:0] s_2060;
  wire [4:0] s_2061;
  wire [4:0] s_2062;
  wire [4:0] s_2063;
  wire [12:0] s_2064;
  wire [12:0] s_2065;
  wire [12:0] s_2066;
  wire [12:0] s_2067;
  wire [12:0] s_2068;
  wire [12:0] s_2069;
  wire [0:0] s_2070;
  wire [12:0] s_2071;
  wire [12:0] s_2072;
  wire [0:0] s_2073;
  wire [0:0] s_2074;
  wire [0:0] s_2075;
  wire [0:0] s_2076;
  wire [0:0] s_2077;
  wire [0:0] s_2078;
  wire [0:0] s_2079;
  wire [0:0] s_2080;
  wire [0:0] s_2081;
  wire [52:0] s_2082;
  wire [0:0] s_2083;
  wire [63:0] s_2084;
  wire [11:0] s_2085;
  wire [0:0] s_2086;
  wire [10:0] s_2087;
  wire [10:0] s_2088;
  wire [12:0] s_2089;
  wire [12:0] s_2090;
  wire [12:0] s_2091;
  wire [12:0] s_2092;
  wire [12:0] s_2093;
  wire [9:0] s_2094;
  wire [51:0] s_2095;
  wire [0:0] s_2096;
  wire [0:0] s_2097;
  wire [10:0] s_2098;
  wire [0:0] s_2099;
  wire [0:0] s_2100;
  wire [0:0] s_2101;
  wire [52:0] s_2102;
  wire [0:0] s_2103;
  wire [0:0] s_2104;
  wire [0:0] s_2105;
  wire [10:0] s_2106;
  wire [0:0] s_2107;
  wire [51:0] s_2108;
  wire [0:0] s_2109;
  wire [0:0] s_2110;
  wire [0:0] s_2111;
  wire [0:0] s_2112;
  wire [10:0] s_2113;
  wire [0:0] s_2114;
  wire [51:0] s_2115;
  wire [0:0] s_2116;
  wire [0:0] s_2117;
  wire [0:0] s_2118;
  wire [0:0] s_2119;

  assign s_0 = s_2109?s_1:s_6;
  dq #(64, 10) dq_s_1 (clk, s_1, s_2);
  assign s_2 = {s_3,s_5};
  assign s_3 = s_4[63];
  assign s_4 = double_sqrt_a;
  assign s_5 = 63'd9221120237041090560;
  assign s_6 = s_2103?s_7:s_10;
  dq #(64, 10) dq_s_7 (clk, s_7, s_8);
  assign s_8 = {s_3,s_9};
  assign s_9 = 63'd9218868437227405312;
  assign s_10 = s_2101?s_11:s_14;
  dq #(64, 10) dq_s_11 (clk, s_11, s_12);
  assign s_12 = {s_3,s_13};
  assign s_13 = 63'd0;
  assign s_14 = s_2096?s_15:s_2084;
  assign s_15 = {s_16,s_19};
  dq #(12, 10) dq_s_16 (clk, s_16, s_17);
  assign s_17 = {s_3,s_18};
  assign s_18 = 11'd0;
  assign s_19 = s_20[51:0];
  dq #(53, 1) dq_s_20 (clk, s_20, s_21);
  assign s_21 = s_2083?s_22:s_2082;
  assign s_22 = s_23[53:1];
  assign s_23 = s_2074?s_24:s_26;
  assign s_24 = s_25 + s_2073;
  assign s_25 = s_26;
  assign s_26 = s_27[53:1];
  dq #(54, 1) dq_s_27 (clk, s_27, s_28);
  assign s_28 = s_29 << s_1349;
  dq #(54, 2) dq_s_29 (clk, s_29, s_30);
  dq #(54, 1) dq_s_30 (clk, s_30, s_31);
  assign s_31 = s_32 >> s_1337;
  dq #(54, 2) dq_s_32 (clk, s_32, s_33);
  assign s_33 = s_34[53:0];
  assign s_34 = s_1330?s_35:s_36;
  assign s_35 = s_36 + s_1329;
  assign s_36 = s_1322?s_37:s_38;
  assign s_37 = s_38 + s_1321;
  assign s_38 = s_1314?s_39:s_40;
  assign s_39 = s_40 + s_1313;
  assign s_40 = s_1306?s_41:s_42;
  assign s_41 = s_42 + s_1305;
  assign s_42 = s_1298?s_43:s_44;
  assign s_43 = s_44 + s_1297;
  assign s_44 = s_1290?s_45:s_46;
  assign s_45 = s_46 + s_1289;
  assign s_46 = s_1282?s_47:s_48;
  assign s_47 = s_48 + s_1281;
  assign s_48 = s_1274?s_49:s_50;
  assign s_49 = s_50 + s_1273;
  assign s_50 = s_1266?s_51:s_52;
  assign s_51 = s_52 + s_1265;
  assign s_52 = s_1258?s_53:s_54;
  assign s_53 = s_54 + s_1257;
  assign s_54 = s_1250?s_55:s_56;
  assign s_55 = s_56 + s_1249;
  assign s_56 = s_1242?s_57:s_58;
  assign s_57 = s_58 + s_1241;
  assign s_58 = s_1234?s_59:s_60;
  assign s_59 = s_60 + s_1233;
  assign s_60 = s_1226?s_61:s_62;
  assign s_61 = s_62 + s_1225;
  assign s_62 = s_1218?s_63:s_64;
  assign s_63 = s_64 + s_1217;
  assign s_64 = s_1210?s_65:s_66;
  assign s_65 = s_66 + s_1209;
  assign s_66 = s_1202?s_67:s_68;
  assign s_67 = s_68 + s_1201;
  assign s_68 = s_1194?s_69:s_70;
  assign s_69 = s_70 + s_1193;
  assign s_70 = s_1186?s_71:s_72;
  assign s_71 = s_72 + s_1185;
  assign s_72 = s_1178?s_73:s_74;
  assign s_73 = s_74 + s_1177;
  assign s_74 = s_1170?s_75:s_76;
  assign s_75 = s_76 + s_1169;
  assign s_76 = s_1162?s_77:s_78;
  assign s_77 = s_78 + s_1161;
  assign s_78 = s_1154?s_79:s_80;
  assign s_79 = s_80 + s_1153;
  assign s_80 = s_1146?s_81:s_82;
  assign s_81 = s_82 + s_1145;
  assign s_82 = s_1138?s_83:s_84;
  assign s_83 = s_84 + s_1137;
  assign s_84 = s_1130?s_85:s_86;
  assign s_85 = s_86 + s_1129;
  assign s_86 = s_1122?s_87:s_88;
  assign s_87 = s_88 + s_1121;
  assign s_88 = s_1114?s_89:s_90;
  assign s_89 = s_90 + s_1113;
  assign s_90 = s_1106?s_91:s_92;
  assign s_91 = s_92 + s_1105;
  assign s_92 = s_1098?s_93:s_94;
  assign s_93 = s_94 + s_1097;
  assign s_94 = s_1090?s_95:s_96;
  assign s_95 = s_96 + s_1089;
  assign s_96 = s_1082?s_97:s_98;
  assign s_97 = s_98 + s_1081;
  assign s_98 = s_1074?s_99:s_100;
  assign s_99 = s_100 + s_1073;
  assign s_100 = s_1066?s_101:s_102;
  assign s_101 = s_102 + s_1065;
  assign s_102 = s_1058?s_103:s_104;
  assign s_103 = s_104 + s_1057;
  assign s_104 = s_1050?s_105:s_106;
  assign s_105 = s_106 + s_1049;
  assign s_106 = s_1042?s_107:s_108;
  assign s_107 = s_108 + s_1041;
  assign s_108 = s_1034?s_109:s_110;
  assign s_109 = s_110 + s_1033;
  assign s_110 = s_1026?s_111:s_112;
  assign s_111 = s_112 + s_1025;
  assign s_112 = s_1018?s_113:s_114;
  assign s_113 = s_114 + s_1017;
  assign s_114 = s_1010?s_115:s_116;
  assign s_115 = s_116 + s_1009;
  assign s_116 = s_1002?s_117:s_118;
  assign s_117 = s_118 + s_1001;
  assign s_118 = s_994?s_119:s_120;
  assign s_119 = s_120 + s_993;
  assign s_120 = s_986?s_121:s_122;
  assign s_121 = s_122 + s_985;
  assign s_122 = s_978?s_123:s_124;
  assign s_123 = s_124 + s_977;
  assign s_124 = s_970?s_125:s_126;
  assign s_125 = s_126 + s_969;
  assign s_126 = s_962?s_127:s_128;
  assign s_127 = s_128 + s_961;
  assign s_128 = s_954?s_129:s_130;
  assign s_129 = s_130 + s_953;
  assign s_130 = s_946?s_131:s_132;
  assign s_131 = s_132 + s_945;
  assign s_132 = s_938?s_133:s_134;
  assign s_133 = s_134 + s_937;
  assign s_134 = s_930?s_135:s_136;
  assign s_135 = s_136 + s_929;
  assign s_136 = s_922?s_137:s_138;
  assign s_137 = s_138 + s_921;
  assign s_138 = s_914?s_139:s_140;
  assign s_139 = s_140 + s_913;
  assign s_140 = s_905?s_141:s_142;
  assign s_141 = s_142 + s_904;
  assign s_142 = s_147?s_143:s_145;
  dq #(109, 3) dq_s_143 (clk, s_143, s_144);
  assign s_144 = s_145 + s_146;
  assign s_145 = 55'd0;
  assign s_146 = 109'd18014398509481984;
  assign s_147 = s_148 <= s_155;
  dq #(110, 3) dq_s_148 (clk, s_148, s_149);
  assign s_149 = s_150 | s_154;
  assign s_150 = s_151 + s_152;
  assign s_151 = 110'd0;
  assign s_152 = s_145 << s_153;
  assign s_153 = 6'd55;
  assign s_154 = 109'd324518553658426726783156020576256;
  assign s_155 = s_156 << s_903;
  assign s_156 = s_899?s_157:s_158;
  assign s_157 = s_158 << s_898;
  assign s_158 = s_159;
  dq #(53, 1) dq_s_159 (clk, s_159, s_160);
  assign s_160 = s_161 << s_172;
  dq #(53, 2) dq_s_161 (clk, s_161, s_162);
  assign s_162 = {s_163,s_171};
  assign s_163 = s_166?s_164:s_165;
  assign s_164 = 1'd0;
  assign s_165 = 1'd1;
  assign s_166 = s_167 == s_170;
  assign s_167 = s_168 - s_169;
  assign s_168 = s_4[62:52];
  assign s_169 = 10'd1023;
  assign s_170 = -11'd1023;
  assign s_171 = s_4[51:0];
  dq #(13, 1) dq_s_172 (clk, s_172, s_173);
  assign s_173 = s_895?s_174:s_889;
  dq #(7, 1) dq_s_174 (clk, s_174, s_175);
  assign s_175 = {s_176,s_883};
  assign s_176 = s_177 & s_541;
  assign s_177 = s_178[5];
  assign s_178 = {s_179,s_535};
  assign s_179 = s_180 & s_369;
  assign s_180 = s_181[4];
  assign s_181 = {s_182,s_363};
  assign s_182 = s_183 & s_285;
  assign s_183 = s_184[3];
  assign s_184 = {s_185,s_279};
  assign s_185 = s_186 & s_245;
  assign s_186 = s_187[2];
  assign s_187 = {s_188,s_239};
  assign s_188 = s_189 & s_227;
  assign s_189 = s_190[1];
  assign s_190 = {s_191,s_223};
  assign s_191 = s_192 & s_221;
  assign s_192 = ~s_193;
  assign s_193 = s_194[1];
  assign s_194 = s_195[3:2];
  assign s_195 = s_196[7:4];
  assign s_196 = s_197[15:8];
  assign s_197 = s_198[31:16];
  assign s_198 = s_199[63:32];
  assign s_199 = {s_200,s_220};
  assign s_200 = {s_201,s_219};
  assign s_201 = {s_202,s_218};
  assign s_202 = {s_203,s_217};
  assign s_203 = {s_204,s_216};
  assign s_204 = {s_205,s_215};
  assign s_205 = {s_206,s_214};
  assign s_206 = {s_207,s_213};
  assign s_207 = {s_208,s_212};
  assign s_208 = {s_209,s_211};
  assign s_209 = {s_162,s_210};
  assign s_210 = 1'd1;
  assign s_211 = 1'd1;
  assign s_212 = 1'd1;
  assign s_213 = 1'd1;
  assign s_214 = 1'd1;
  assign s_215 = 1'd1;
  assign s_216 = 1'd1;
  assign s_217 = 1'd1;
  assign s_218 = 1'd1;
  assign s_219 = 1'd1;
  assign s_220 = 1'd1;
  assign s_221 = ~s_222;
  assign s_222 = s_194[0];
  assign s_223 = s_224 & s_226;
  assign s_224 = ~s_225;
  assign s_225 = s_194[1];
  assign s_226 = s_194[0];
  assign s_227 = s_228[1];
  assign s_228 = {s_229,s_235};
  assign s_229 = s_230 & s_233;
  assign s_230 = ~s_231;
  assign s_231 = s_232[1];
  assign s_232 = s_195[1:0];
  assign s_233 = ~s_234;
  assign s_234 = s_232[0];
  assign s_235 = s_236 & s_238;
  assign s_236 = ~s_237;
  assign s_237 = s_232[1];
  assign s_238 = s_232[0];
  assign s_239 = {s_240,s_242};
  assign s_240 = s_189 & s_241;
  assign s_241 = ~s_227;
  assign s_242 = s_189?s_243:s_244;
  assign s_243 = s_228[0:0];
  assign s_244 = s_190[0:0];
  assign s_245 = s_246[2];
  assign s_246 = {s_247,s_273};
  assign s_247 = s_248 & s_261;
  assign s_248 = s_249[1];
  assign s_249 = {s_250,s_257};
  assign s_250 = s_251 & s_255;
  assign s_251 = ~s_252;
  assign s_252 = s_253[1];
  assign s_253 = s_254[3:2];
  assign s_254 = s_196[3:0];
  assign s_255 = ~s_256;
  assign s_256 = s_253[0];
  assign s_257 = s_258 & s_260;
  assign s_258 = ~s_259;
  assign s_259 = s_253[1];
  assign s_260 = s_253[0];
  assign s_261 = s_262[1];
  assign s_262 = {s_263,s_269};
  assign s_263 = s_264 & s_267;
  assign s_264 = ~s_265;
  assign s_265 = s_266[1];
  assign s_266 = s_254[1:0];
  assign s_267 = ~s_268;
  assign s_268 = s_266[0];
  assign s_269 = s_270 & s_272;
  assign s_270 = ~s_271;
  assign s_271 = s_266[1];
  assign s_272 = s_266[0];
  assign s_273 = {s_274,s_276};
  assign s_274 = s_248 & s_275;
  assign s_275 = ~s_261;
  assign s_276 = s_248?s_277:s_278;
  assign s_277 = s_262[0:0];
  assign s_278 = s_249[0:0];
  assign s_279 = {s_280,s_282};
  assign s_280 = s_186 & s_281;
  assign s_281 = ~s_245;
  assign s_282 = s_186?s_283:s_284;
  assign s_283 = s_246[1:0];
  assign s_284 = s_187[1:0];
  assign s_285 = s_286[3];
  assign s_286 = {s_287,s_357};
  assign s_287 = s_288 & s_323;
  assign s_288 = s_289[2];
  assign s_289 = {s_290,s_317};
  assign s_290 = s_291 & s_305;
  assign s_291 = s_292[1];
  assign s_292 = {s_293,s_301};
  assign s_293 = s_294 & s_299;
  assign s_294 = ~s_295;
  assign s_295 = s_296[1];
  assign s_296 = s_297[3:2];
  assign s_297 = s_298[7:4];
  assign s_298 = s_197[7:0];
  assign s_299 = ~s_300;
  assign s_300 = s_296[0];
  assign s_301 = s_302 & s_304;
  assign s_302 = ~s_303;
  assign s_303 = s_296[1];
  assign s_304 = s_296[0];
  assign s_305 = s_306[1];
  assign s_306 = {s_307,s_313};
  assign s_307 = s_308 & s_311;
  assign s_308 = ~s_309;
  assign s_309 = s_310[1];
  assign s_310 = s_297[1:0];
  assign s_311 = ~s_312;
  assign s_312 = s_310[0];
  assign s_313 = s_314 & s_316;
  assign s_314 = ~s_315;
  assign s_315 = s_310[1];
  assign s_316 = s_310[0];
  assign s_317 = {s_318,s_320};
  assign s_318 = s_291 & s_319;
  assign s_319 = ~s_305;
  assign s_320 = s_291?s_321:s_322;
  assign s_321 = s_306[0:0];
  assign s_322 = s_292[0:0];
  assign s_323 = s_324[2];
  assign s_324 = {s_325,s_351};
  assign s_325 = s_326 & s_339;
  assign s_326 = s_327[1];
  assign s_327 = {s_328,s_335};
  assign s_328 = s_329 & s_333;
  assign s_329 = ~s_330;
  assign s_330 = s_331[1];
  assign s_331 = s_332[3:2];
  assign s_332 = s_298[3:0];
  assign s_333 = ~s_334;
  assign s_334 = s_331[0];
  assign s_335 = s_336 & s_338;
  assign s_336 = ~s_337;
  assign s_337 = s_331[1];
  assign s_338 = s_331[0];
  assign s_339 = s_340[1];
  assign s_340 = {s_341,s_347};
  assign s_341 = s_342 & s_345;
  assign s_342 = ~s_343;
  assign s_343 = s_344[1];
  assign s_344 = s_332[1:0];
  assign s_345 = ~s_346;
  assign s_346 = s_344[0];
  assign s_347 = s_348 & s_350;
  assign s_348 = ~s_349;
  assign s_349 = s_344[1];
  assign s_350 = s_344[0];
  assign s_351 = {s_352,s_354};
  assign s_352 = s_326 & s_353;
  assign s_353 = ~s_339;
  assign s_354 = s_326?s_355:s_356;
  assign s_355 = s_340[0:0];
  assign s_356 = s_327[0:0];
  assign s_357 = {s_358,s_360};
  assign s_358 = s_288 & s_359;
  assign s_359 = ~s_323;
  assign s_360 = s_288?s_361:s_362;
  assign s_361 = s_324[1:0];
  assign s_362 = s_289[1:0];
  assign s_363 = {s_364,s_366};
  assign s_364 = s_183 & s_365;
  assign s_365 = ~s_285;
  assign s_366 = s_183?s_367:s_368;
  assign s_367 = s_286[2:0];
  assign s_368 = s_184[2:0];
  assign s_369 = s_370[4];
  assign s_370 = {s_371,s_529};
  assign s_371 = s_372 & s_451;
  assign s_372 = s_373[3];
  assign s_373 = {s_374,s_445};
  assign s_374 = s_375 & s_411;
  assign s_375 = s_376[2];
  assign s_376 = {s_377,s_405};
  assign s_377 = s_378 & s_393;
  assign s_378 = s_379[1];
  assign s_379 = {s_380,s_389};
  assign s_380 = s_381 & s_387;
  assign s_381 = ~s_382;
  assign s_382 = s_383[1];
  assign s_383 = s_384[3:2];
  assign s_384 = s_385[7:4];
  assign s_385 = s_386[15:8];
  assign s_386 = s_198[15:0];
  assign s_387 = ~s_388;
  assign s_388 = s_383[0];
  assign s_389 = s_390 & s_392;
  assign s_390 = ~s_391;
  assign s_391 = s_383[1];
  assign s_392 = s_383[0];
  assign s_393 = s_394[1];
  assign s_394 = {s_395,s_401};
  assign s_395 = s_396 & s_399;
  assign s_396 = ~s_397;
  assign s_397 = s_398[1];
  assign s_398 = s_384[1:0];
  assign s_399 = ~s_400;
  assign s_400 = s_398[0];
  assign s_401 = s_402 & s_404;
  assign s_402 = ~s_403;
  assign s_403 = s_398[1];
  assign s_404 = s_398[0];
  assign s_405 = {s_406,s_408};
  assign s_406 = s_378 & s_407;
  assign s_407 = ~s_393;
  assign s_408 = s_378?s_409:s_410;
  assign s_409 = s_394[0:0];
  assign s_410 = s_379[0:0];
  assign s_411 = s_412[2];
  assign s_412 = {s_413,s_439};
  assign s_413 = s_414 & s_427;
  assign s_414 = s_415[1];
  assign s_415 = {s_416,s_423};
  assign s_416 = s_417 & s_421;
  assign s_417 = ~s_418;
  assign s_418 = s_419[1];
  assign s_419 = s_420[3:2];
  assign s_420 = s_385[3:0];
  assign s_421 = ~s_422;
  assign s_422 = s_419[0];
  assign s_423 = s_424 & s_426;
  assign s_424 = ~s_425;
  assign s_425 = s_419[1];
  assign s_426 = s_419[0];
  assign s_427 = s_428[1];
  assign s_428 = {s_429,s_435};
  assign s_429 = s_430 & s_433;
  assign s_430 = ~s_431;
  assign s_431 = s_432[1];
  assign s_432 = s_420[1:0];
  assign s_433 = ~s_434;
  assign s_434 = s_432[0];
  assign s_435 = s_436 & s_438;
  assign s_436 = ~s_437;
  assign s_437 = s_432[1];
  assign s_438 = s_432[0];
  assign s_439 = {s_440,s_442};
  assign s_440 = s_414 & s_441;
  assign s_441 = ~s_427;
  assign s_442 = s_414?s_443:s_444;
  assign s_443 = s_428[0:0];
  assign s_444 = s_415[0:0];
  assign s_445 = {s_446,s_448};
  assign s_446 = s_375 & s_447;
  assign s_447 = ~s_411;
  assign s_448 = s_375?s_449:s_450;
  assign s_449 = s_412[1:0];
  assign s_450 = s_376[1:0];
  assign s_451 = s_452[3];
  assign s_452 = {s_453,s_523};
  assign s_453 = s_454 & s_489;
  assign s_454 = s_455[2];
  assign s_455 = {s_456,s_483};
  assign s_456 = s_457 & s_471;
  assign s_457 = s_458[1];
  assign s_458 = {s_459,s_467};
  assign s_459 = s_460 & s_465;
  assign s_460 = ~s_461;
  assign s_461 = s_462[1];
  assign s_462 = s_463[3:2];
  assign s_463 = s_464[7:4];
  assign s_464 = s_386[7:0];
  assign s_465 = ~s_466;
  assign s_466 = s_462[0];
  assign s_467 = s_468 & s_470;
  assign s_468 = ~s_469;
  assign s_469 = s_462[1];
  assign s_470 = s_462[0];
  assign s_471 = s_472[1];
  assign s_472 = {s_473,s_479};
  assign s_473 = s_474 & s_477;
  assign s_474 = ~s_475;
  assign s_475 = s_476[1];
  assign s_476 = s_463[1:0];
  assign s_477 = ~s_478;
  assign s_478 = s_476[0];
  assign s_479 = s_480 & s_482;
  assign s_480 = ~s_481;
  assign s_481 = s_476[1];
  assign s_482 = s_476[0];
  assign s_483 = {s_484,s_486};
  assign s_484 = s_457 & s_485;
  assign s_485 = ~s_471;
  assign s_486 = s_457?s_487:s_488;
  assign s_487 = s_472[0:0];
  assign s_488 = s_458[0:0];
  assign s_489 = s_490[2];
  assign s_490 = {s_491,s_517};
  assign s_491 = s_492 & s_505;
  assign s_492 = s_493[1];
  assign s_493 = {s_494,s_501};
  assign s_494 = s_495 & s_499;
  assign s_495 = ~s_496;
  assign s_496 = s_497[1];
  assign s_497 = s_498[3:2];
  assign s_498 = s_464[3:0];
  assign s_499 = ~s_500;
  assign s_500 = s_497[0];
  assign s_501 = s_502 & s_504;
  assign s_502 = ~s_503;
  assign s_503 = s_497[1];
  assign s_504 = s_497[0];
  assign s_505 = s_506[1];
  assign s_506 = {s_507,s_513};
  assign s_507 = s_508 & s_511;
  assign s_508 = ~s_509;
  assign s_509 = s_510[1];
  assign s_510 = s_498[1:0];
  assign s_511 = ~s_512;
  assign s_512 = s_510[0];
  assign s_513 = s_514 & s_516;
  assign s_514 = ~s_515;
  assign s_515 = s_510[1];
  assign s_516 = s_510[0];
  assign s_517 = {s_518,s_520};
  assign s_518 = s_492 & s_519;
  assign s_519 = ~s_505;
  assign s_520 = s_492?s_521:s_522;
  assign s_521 = s_506[0:0];
  assign s_522 = s_493[0:0];
  assign s_523 = {s_524,s_526};
  assign s_524 = s_454 & s_525;
  assign s_525 = ~s_489;
  assign s_526 = s_454?s_527:s_528;
  assign s_527 = s_490[1:0];
  assign s_528 = s_455[1:0];
  assign s_529 = {s_530,s_532};
  assign s_530 = s_372 & s_531;
  assign s_531 = ~s_451;
  assign s_532 = s_372?s_533:s_534;
  assign s_533 = s_452[2:0];
  assign s_534 = s_373[2:0];
  assign s_535 = {s_536,s_538};
  assign s_536 = s_180 & s_537;
  assign s_537 = ~s_369;
  assign s_538 = s_180?s_539:s_540;
  assign s_539 = s_370[3:0];
  assign s_540 = s_181[3:0];
  assign s_541 = s_542[5];
  assign s_542 = {s_543,s_877};
  assign s_543 = s_544 & s_711;
  assign s_544 = s_545[4];
  assign s_545 = {s_546,s_705};
  assign s_546 = s_547 & s_627;
  assign s_547 = s_548[3];
  assign s_548 = {s_549,s_621};
  assign s_549 = s_550 & s_587;
  assign s_550 = s_551[2];
  assign s_551 = {s_552,s_581};
  assign s_552 = s_553 & s_569;
  assign s_553 = s_554[1];
  assign s_554 = {s_555,s_565};
  assign s_555 = s_556 & s_563;
  assign s_556 = ~s_557;
  assign s_557 = s_558[1];
  assign s_558 = s_559[3:2];
  assign s_559 = s_560[7:4];
  assign s_560 = s_561[15:8];
  assign s_561 = s_562[31:16];
  assign s_562 = s_199[31:0];
  assign s_563 = ~s_564;
  assign s_564 = s_558[0];
  assign s_565 = s_566 & s_568;
  assign s_566 = ~s_567;
  assign s_567 = s_558[1];
  assign s_568 = s_558[0];
  assign s_569 = s_570[1];
  assign s_570 = {s_571,s_577};
  assign s_571 = s_572 & s_575;
  assign s_572 = ~s_573;
  assign s_573 = s_574[1];
  assign s_574 = s_559[1:0];
  assign s_575 = ~s_576;
  assign s_576 = s_574[0];
  assign s_577 = s_578 & s_580;
  assign s_578 = ~s_579;
  assign s_579 = s_574[1];
  assign s_580 = s_574[0];
  assign s_581 = {s_582,s_584};
  assign s_582 = s_553 & s_583;
  assign s_583 = ~s_569;
  assign s_584 = s_553?s_585:s_586;
  assign s_585 = s_570[0:0];
  assign s_586 = s_554[0:0];
  assign s_587 = s_588[2];
  assign s_588 = {s_589,s_615};
  assign s_589 = s_590 & s_603;
  assign s_590 = s_591[1];
  assign s_591 = {s_592,s_599};
  assign s_592 = s_593 & s_597;
  assign s_593 = ~s_594;
  assign s_594 = s_595[1];
  assign s_595 = s_596[3:2];
  assign s_596 = s_560[3:0];
  assign s_597 = ~s_598;
  assign s_598 = s_595[0];
  assign s_599 = s_600 & s_602;
  assign s_600 = ~s_601;
  assign s_601 = s_595[1];
  assign s_602 = s_595[0];
  assign s_603 = s_604[1];
  assign s_604 = {s_605,s_611};
  assign s_605 = s_606 & s_609;
  assign s_606 = ~s_607;
  assign s_607 = s_608[1];
  assign s_608 = s_596[1:0];
  assign s_609 = ~s_610;
  assign s_610 = s_608[0];
  assign s_611 = s_612 & s_614;
  assign s_612 = ~s_613;
  assign s_613 = s_608[1];
  assign s_614 = s_608[0];
  assign s_615 = {s_616,s_618};
  assign s_616 = s_590 & s_617;
  assign s_617 = ~s_603;
  assign s_618 = s_590?s_619:s_620;
  assign s_619 = s_604[0:0];
  assign s_620 = s_591[0:0];
  assign s_621 = {s_622,s_624};
  assign s_622 = s_550 & s_623;
  assign s_623 = ~s_587;
  assign s_624 = s_550?s_625:s_626;
  assign s_625 = s_588[1:0];
  assign s_626 = s_551[1:0];
  assign s_627 = s_628[3];
  assign s_628 = {s_629,s_699};
  assign s_629 = s_630 & s_665;
  assign s_630 = s_631[2];
  assign s_631 = {s_632,s_659};
  assign s_632 = s_633 & s_647;
  assign s_633 = s_634[1];
  assign s_634 = {s_635,s_643};
  assign s_635 = s_636 & s_641;
  assign s_636 = ~s_637;
  assign s_637 = s_638[1];
  assign s_638 = s_639[3:2];
  assign s_639 = s_640[7:4];
  assign s_640 = s_561[7:0];
  assign s_641 = ~s_642;
  assign s_642 = s_638[0];
  assign s_643 = s_644 & s_646;
  assign s_644 = ~s_645;
  assign s_645 = s_638[1];
  assign s_646 = s_638[0];
  assign s_647 = s_648[1];
  assign s_648 = {s_649,s_655};
  assign s_649 = s_650 & s_653;
  assign s_650 = ~s_651;
  assign s_651 = s_652[1];
  assign s_652 = s_639[1:0];
  assign s_653 = ~s_654;
  assign s_654 = s_652[0];
  assign s_655 = s_656 & s_658;
  assign s_656 = ~s_657;
  assign s_657 = s_652[1];
  assign s_658 = s_652[0];
  assign s_659 = {s_660,s_662};
  assign s_660 = s_633 & s_661;
  assign s_661 = ~s_647;
  assign s_662 = s_633?s_663:s_664;
  assign s_663 = s_648[0:0];
  assign s_664 = s_634[0:0];
  assign s_665 = s_666[2];
  assign s_666 = {s_667,s_693};
  assign s_667 = s_668 & s_681;
  assign s_668 = s_669[1];
  assign s_669 = {s_670,s_677};
  assign s_670 = s_671 & s_675;
  assign s_671 = ~s_672;
  assign s_672 = s_673[1];
  assign s_673 = s_674[3:2];
  assign s_674 = s_640[3:0];
  assign s_675 = ~s_676;
  assign s_676 = s_673[0];
  assign s_677 = s_678 & s_680;
  assign s_678 = ~s_679;
  assign s_679 = s_673[1];
  assign s_680 = s_673[0];
  assign s_681 = s_682[1];
  assign s_682 = {s_683,s_689};
  assign s_683 = s_684 & s_687;
  assign s_684 = ~s_685;
  assign s_685 = s_686[1];
  assign s_686 = s_674[1:0];
  assign s_687 = ~s_688;
  assign s_688 = s_686[0];
  assign s_689 = s_690 & s_692;
  assign s_690 = ~s_691;
  assign s_691 = s_686[1];
  assign s_692 = s_686[0];
  assign s_693 = {s_694,s_696};
  assign s_694 = s_668 & s_695;
  assign s_695 = ~s_681;
  assign s_696 = s_668?s_697:s_698;
  assign s_697 = s_682[0:0];
  assign s_698 = s_669[0:0];
  assign s_699 = {s_700,s_702};
  assign s_700 = s_630 & s_701;
  assign s_701 = ~s_665;
  assign s_702 = s_630?s_703:s_704;
  assign s_703 = s_666[1:0];
  assign s_704 = s_631[1:0];
  assign s_705 = {s_706,s_708};
  assign s_706 = s_547 & s_707;
  assign s_707 = ~s_627;
  assign s_708 = s_547?s_709:s_710;
  assign s_709 = s_628[2:0];
  assign s_710 = s_548[2:0];
  assign s_711 = s_712[4];
  assign s_712 = {s_713,s_871};
  assign s_713 = s_714 & s_793;
  assign s_714 = s_715[3];
  assign s_715 = {s_716,s_787};
  assign s_716 = s_717 & s_753;
  assign s_717 = s_718[2];
  assign s_718 = {s_719,s_747};
  assign s_719 = s_720 & s_735;
  assign s_720 = s_721[1];
  assign s_721 = {s_722,s_731};
  assign s_722 = s_723 & s_729;
  assign s_723 = ~s_724;
  assign s_724 = s_725[1];
  assign s_725 = s_726[3:2];
  assign s_726 = s_727[7:4];
  assign s_727 = s_728[15:8];
  assign s_728 = s_562[15:0];
  assign s_729 = ~s_730;
  assign s_730 = s_725[0];
  assign s_731 = s_732 & s_734;
  assign s_732 = ~s_733;
  assign s_733 = s_725[1];
  assign s_734 = s_725[0];
  assign s_735 = s_736[1];
  assign s_736 = {s_737,s_743};
  assign s_737 = s_738 & s_741;
  assign s_738 = ~s_739;
  assign s_739 = s_740[1];
  assign s_740 = s_726[1:0];
  assign s_741 = ~s_742;
  assign s_742 = s_740[0];
  assign s_743 = s_744 & s_746;
  assign s_744 = ~s_745;
  assign s_745 = s_740[1];
  assign s_746 = s_740[0];
  assign s_747 = {s_748,s_750};
  assign s_748 = s_720 & s_749;
  assign s_749 = ~s_735;
  assign s_750 = s_720?s_751:s_752;
  assign s_751 = s_736[0:0];
  assign s_752 = s_721[0:0];
  assign s_753 = s_754[2];
  assign s_754 = {s_755,s_781};
  assign s_755 = s_756 & s_769;
  assign s_756 = s_757[1];
  assign s_757 = {s_758,s_765};
  assign s_758 = s_759 & s_763;
  assign s_759 = ~s_760;
  assign s_760 = s_761[1];
  assign s_761 = s_762[3:2];
  assign s_762 = s_727[3:0];
  assign s_763 = ~s_764;
  assign s_764 = s_761[0];
  assign s_765 = s_766 & s_768;
  assign s_766 = ~s_767;
  assign s_767 = s_761[1];
  assign s_768 = s_761[0];
  assign s_769 = s_770[1];
  assign s_770 = {s_771,s_777};
  assign s_771 = s_772 & s_775;
  assign s_772 = ~s_773;
  assign s_773 = s_774[1];
  assign s_774 = s_762[1:0];
  assign s_775 = ~s_776;
  assign s_776 = s_774[0];
  assign s_777 = s_778 & s_780;
  assign s_778 = ~s_779;
  assign s_779 = s_774[1];
  assign s_780 = s_774[0];
  assign s_781 = {s_782,s_784};
  assign s_782 = s_756 & s_783;
  assign s_783 = ~s_769;
  assign s_784 = s_756?s_785:s_786;
  assign s_785 = s_770[0:0];
  assign s_786 = s_757[0:0];
  assign s_787 = {s_788,s_790};
  assign s_788 = s_717 & s_789;
  assign s_789 = ~s_753;
  assign s_790 = s_717?s_791:s_792;
  assign s_791 = s_754[1:0];
  assign s_792 = s_718[1:0];
  assign s_793 = s_794[3];
  assign s_794 = {s_795,s_865};
  assign s_795 = s_796 & s_831;
  assign s_796 = s_797[2];
  assign s_797 = {s_798,s_825};
  assign s_798 = s_799 & s_813;
  assign s_799 = s_800[1];
  assign s_800 = {s_801,s_809};
  assign s_801 = s_802 & s_807;
  assign s_802 = ~s_803;
  assign s_803 = s_804[1];
  assign s_804 = s_805[3:2];
  assign s_805 = s_806[7:4];
  assign s_806 = s_728[7:0];
  assign s_807 = ~s_808;
  assign s_808 = s_804[0];
  assign s_809 = s_810 & s_812;
  assign s_810 = ~s_811;
  assign s_811 = s_804[1];
  assign s_812 = s_804[0];
  assign s_813 = s_814[1];
  assign s_814 = {s_815,s_821};
  assign s_815 = s_816 & s_819;
  assign s_816 = ~s_817;
  assign s_817 = s_818[1];
  assign s_818 = s_805[1:0];
  assign s_819 = ~s_820;
  assign s_820 = s_818[0];
  assign s_821 = s_822 & s_824;
  assign s_822 = ~s_823;
  assign s_823 = s_818[1];
  assign s_824 = s_818[0];
  assign s_825 = {s_826,s_828};
  assign s_826 = s_799 & s_827;
  assign s_827 = ~s_813;
  assign s_828 = s_799?s_829:s_830;
  assign s_829 = s_814[0:0];
  assign s_830 = s_800[0:0];
  assign s_831 = s_832[2];
  assign s_832 = {s_833,s_859};
  assign s_833 = s_834 & s_847;
  assign s_834 = s_835[1];
  assign s_835 = {s_836,s_843};
  assign s_836 = s_837 & s_841;
  assign s_837 = ~s_838;
  assign s_838 = s_839[1];
  assign s_839 = s_840[3:2];
  assign s_840 = s_806[3:0];
  assign s_841 = ~s_842;
  assign s_842 = s_839[0];
  assign s_843 = s_844 & s_846;
  assign s_844 = ~s_845;
  assign s_845 = s_839[1];
  assign s_846 = s_839[0];
  assign s_847 = s_848[1];
  assign s_848 = {s_849,s_855};
  assign s_849 = s_850 & s_853;
  assign s_850 = ~s_851;
  assign s_851 = s_852[1];
  assign s_852 = s_840[1:0];
  assign s_853 = ~s_854;
  assign s_854 = s_852[0];
  assign s_855 = s_856 & s_858;
  assign s_856 = ~s_857;
  assign s_857 = s_852[1];
  assign s_858 = s_852[0];
  assign s_859 = {s_860,s_862};
  assign s_860 = s_834 & s_861;
  assign s_861 = ~s_847;
  assign s_862 = s_834?s_863:s_864;
  assign s_863 = s_848[0:0];
  assign s_864 = s_835[0:0];
  assign s_865 = {s_866,s_868};
  assign s_866 = s_796 & s_867;
  assign s_867 = ~s_831;
  assign s_868 = s_796?s_869:s_870;
  assign s_869 = s_832[1:0];
  assign s_870 = s_797[1:0];
  assign s_871 = {s_872,s_874};
  assign s_872 = s_714 & s_873;
  assign s_873 = ~s_793;
  assign s_874 = s_714?s_875:s_876;
  assign s_875 = s_794[2:0];
  assign s_876 = s_715[2:0];
  assign s_877 = {s_878,s_880};
  assign s_878 = s_544 & s_879;
  assign s_879 = ~s_711;
  assign s_880 = s_544?s_881:s_882;
  assign s_881 = s_712[3:0];
  assign s_882 = s_545[3:0];
  assign s_883 = {s_884,s_886};
  assign s_884 = s_177 & s_885;
  assign s_885 = ~s_541;
  assign s_886 = s_177?s_887:s_888;
  assign s_887 = s_542[4:0];
  assign s_888 = s_178[4:0];
  dq #(13, 1) dq_s_889 (clk, s_889, s_890);
  assign s_890 = s_891 - s_894;
  assign s_891 = $signed(s_892);
  assign s_892 = s_166?s_893:s_167;
  assign s_893 = -11'd1022;
  assign s_894 = -13'd2044;
  assign s_895 = s_896 <= s_897;
  assign s_896 = s_174;
  dq #(13, 1) dq_s_897 (clk, s_897, s_890);
  assign s_898 = 1'd1;
  assign s_899 = s_900[0];
  dq #(13, 1) dq_s_900 (clk, s_900, s_901);
  assign s_901 = s_902 - s_172;
  dq #(13, 2) dq_s_902 (clk, s_902, s_891);
  assign s_903 = 6'd54;
  assign s_904 = 109'd9007199254740992;
  assign s_905 = s_906 <= s_155;
  assign s_906 = s_907 | s_912;
  assign s_907 = s_908 + s_910;
  assign s_908 = s_147?s_909:s_151;
  dq #(110, 3) dq_s_909 (clk, s_909, s_149);
  assign s_910 = s_142 << s_911;
  assign s_911 = 6'd54;
  assign s_912 = 107'd81129638414606681695789005144064;
  assign s_913 = 109'd4503599627370496;
  assign s_914 = s_915 <= s_155;
  assign s_915 = s_916 | s_920;
  assign s_916 = s_917 + s_918;
  assign s_917 = s_905?s_906:s_908;
  assign s_918 = s_140 << s_919;
  assign s_919 = 6'd53;
  assign s_920 = 105'd20282409603651670423947251286016;
  assign s_921 = 109'd2251799813685248;
  assign s_922 = s_923 <= s_155;
  assign s_923 = s_924 | s_928;
  assign s_924 = s_925 + s_926;
  assign s_925 = s_914?s_915:s_917;
  assign s_926 = s_138 << s_927;
  assign s_927 = 6'd52;
  assign s_928 = 103'd5070602400912917605986812821504;
  assign s_929 = 109'd1125899906842624;
  assign s_930 = s_931 <= s_155;
  assign s_931 = s_932 | s_936;
  assign s_932 = s_933 + s_934;
  assign s_933 = s_922?s_923:s_925;
  assign s_934 = s_136 << s_935;
  assign s_935 = 6'd51;
  assign s_936 = 101'd1267650600228229401496703205376;
  assign s_937 = 109'd562949953421312;
  assign s_938 = s_939 <= s_155;
  assign s_939 = s_940 | s_944;
  assign s_940 = s_941 + s_942;
  assign s_941 = s_930?s_931:s_933;
  assign s_942 = s_134 << s_943;
  assign s_943 = 6'd50;
  assign s_944 = 99'd316912650057057350374175801344;
  assign s_945 = 109'd281474976710656;
  assign s_946 = s_947 <= s_155;
  assign s_947 = s_948 | s_952;
  assign s_948 = s_949 + s_950;
  assign s_949 = s_938?s_939:s_941;
  assign s_950 = s_132 << s_951;
  assign s_951 = 6'd49;
  assign s_952 = 97'd79228162514264337593543950336;
  assign s_953 = 109'd140737488355328;
  assign s_954 = s_955 <= s_155;
  assign s_955 = s_956 | s_960;
  assign s_956 = s_957 + s_958;
  assign s_957 = s_946?s_947:s_949;
  assign s_958 = s_130 << s_959;
  assign s_959 = 6'd48;
  assign s_960 = 95'd19807040628566084398385987584;
  assign s_961 = 109'd70368744177664;
  assign s_962 = s_963 <= s_155;
  assign s_963 = s_964 | s_968;
  assign s_964 = s_965 + s_966;
  assign s_965 = s_954?s_955:s_957;
  assign s_966 = s_128 << s_967;
  assign s_967 = 6'd47;
  assign s_968 = 93'd4951760157141521099596496896;
  assign s_969 = 109'd35184372088832;
  assign s_970 = s_971 <= s_155;
  assign s_971 = s_972 | s_976;
  assign s_972 = s_973 + s_974;
  assign s_973 = s_962?s_963:s_965;
  assign s_974 = s_126 << s_975;
  assign s_975 = 6'd46;
  assign s_976 = 91'd1237940039285380274899124224;
  assign s_977 = 109'd17592186044416;
  assign s_978 = s_979 <= s_155;
  assign s_979 = s_980 | s_984;
  assign s_980 = s_981 + s_982;
  assign s_981 = s_970?s_971:s_973;
  assign s_982 = s_124 << s_983;
  assign s_983 = 6'd45;
  assign s_984 = 89'd309485009821345068724781056;
  assign s_985 = 109'd8796093022208;
  assign s_986 = s_987 <= s_155;
  assign s_987 = s_988 | s_992;
  assign s_988 = s_989 + s_990;
  assign s_989 = s_978?s_979:s_981;
  assign s_990 = s_122 << s_991;
  assign s_991 = 6'd44;
  assign s_992 = 87'd77371252455336267181195264;
  assign s_993 = 109'd4398046511104;
  assign s_994 = s_995 <= s_155;
  assign s_995 = s_996 | s_1000;
  assign s_996 = s_997 + s_998;
  assign s_997 = s_986?s_987:s_989;
  assign s_998 = s_120 << s_999;
  assign s_999 = 6'd43;
  assign s_1000 = 85'd19342813113834066795298816;
  assign s_1001 = 109'd2199023255552;
  assign s_1002 = s_1003 <= s_155;
  assign s_1003 = s_1004 | s_1008;
  assign s_1004 = s_1005 + s_1006;
  assign s_1005 = s_994?s_995:s_997;
  assign s_1006 = s_118 << s_1007;
  assign s_1007 = 6'd42;
  assign s_1008 = 83'd4835703278458516698824704;
  assign s_1009 = 109'd1099511627776;
  assign s_1010 = s_1011 <= s_155;
  assign s_1011 = s_1012 | s_1016;
  assign s_1012 = s_1013 + s_1014;
  assign s_1013 = s_1002?s_1003:s_1005;
  assign s_1014 = s_116 << s_1015;
  assign s_1015 = 6'd41;
  assign s_1016 = 81'd1208925819614629174706176;
  assign s_1017 = 109'd549755813888;
  assign s_1018 = s_1019 <= s_155;
  assign s_1019 = s_1020 | s_1024;
  assign s_1020 = s_1021 + s_1022;
  assign s_1021 = s_1010?s_1011:s_1013;
  assign s_1022 = s_114 << s_1023;
  assign s_1023 = 6'd40;
  assign s_1024 = 79'd302231454903657293676544;
  assign s_1025 = 109'd274877906944;
  assign s_1026 = s_1027 <= s_155;
  assign s_1027 = s_1028 | s_1032;
  assign s_1028 = s_1029 + s_1030;
  assign s_1029 = s_1018?s_1019:s_1021;
  assign s_1030 = s_112 << s_1031;
  assign s_1031 = 6'd39;
  assign s_1032 = 77'd75557863725914323419136;
  assign s_1033 = 109'd137438953472;
  assign s_1034 = s_1035 <= s_155;
  assign s_1035 = s_1036 | s_1040;
  assign s_1036 = s_1037 + s_1038;
  assign s_1037 = s_1026?s_1027:s_1029;
  assign s_1038 = s_110 << s_1039;
  assign s_1039 = 6'd38;
  assign s_1040 = 75'd18889465931478580854784;
  assign s_1041 = 109'd68719476736;
  assign s_1042 = s_1043 <= s_155;
  assign s_1043 = s_1044 | s_1048;
  assign s_1044 = s_1045 + s_1046;
  assign s_1045 = s_1034?s_1035:s_1037;
  assign s_1046 = s_108 << s_1047;
  assign s_1047 = 6'd37;
  assign s_1048 = 73'd4722366482869645213696;
  assign s_1049 = 109'd34359738368;
  assign s_1050 = s_1051 <= s_155;
  assign s_1051 = s_1052 | s_1056;
  assign s_1052 = s_1053 + s_1054;
  assign s_1053 = s_1042?s_1043:s_1045;
  assign s_1054 = s_106 << s_1055;
  assign s_1055 = 6'd36;
  assign s_1056 = 71'd1180591620717411303424;
  assign s_1057 = 109'd17179869184;
  assign s_1058 = s_1059 <= s_155;
  assign s_1059 = s_1060 | s_1064;
  assign s_1060 = s_1061 + s_1062;
  assign s_1061 = s_1050?s_1051:s_1053;
  assign s_1062 = s_104 << s_1063;
  assign s_1063 = 6'd35;
  assign s_1064 = 69'd295147905179352825856;
  assign s_1065 = 109'd8589934592;
  assign s_1066 = s_1067 <= s_155;
  assign s_1067 = s_1068 | s_1072;
  assign s_1068 = s_1069 + s_1070;
  assign s_1069 = s_1058?s_1059:s_1061;
  assign s_1070 = s_102 << s_1071;
  assign s_1071 = 6'd34;
  assign s_1072 = 67'd73786976294838206464;
  assign s_1073 = 109'd4294967296;
  assign s_1074 = s_1075 <= s_155;
  assign s_1075 = s_1076 | s_1080;
  assign s_1076 = s_1077 + s_1078;
  assign s_1077 = s_1066?s_1067:s_1069;
  assign s_1078 = s_100 << s_1079;
  assign s_1079 = 6'd33;
  assign s_1080 = 65'd18446744073709551616;
  assign s_1081 = 109'd2147483648;
  assign s_1082 = s_1083 <= s_155;
  assign s_1083 = s_1084 | s_1088;
  assign s_1084 = s_1085 + s_1086;
  assign s_1085 = s_1074?s_1075:s_1077;
  assign s_1086 = s_98 << s_1087;
  assign s_1087 = 6'd32;
  assign s_1088 = 63'd4611686018427387904;
  assign s_1089 = 109'd1073741824;
  assign s_1090 = s_1091 <= s_155;
  assign s_1091 = s_1092 | s_1096;
  assign s_1092 = s_1093 + s_1094;
  assign s_1093 = s_1082?s_1083:s_1085;
  assign s_1094 = s_96 << s_1095;
  assign s_1095 = 5'd31;
  assign s_1096 = 61'd1152921504606846976;
  assign s_1097 = 109'd536870912;
  assign s_1098 = s_1099 <= s_155;
  assign s_1099 = s_1100 | s_1104;
  assign s_1100 = s_1101 + s_1102;
  assign s_1101 = s_1090?s_1091:s_1093;
  assign s_1102 = s_94 << s_1103;
  assign s_1103 = 5'd30;
  assign s_1104 = 59'd288230376151711744;
  assign s_1105 = 109'd268435456;
  assign s_1106 = s_1107 <= s_155;
  assign s_1107 = s_1108 | s_1112;
  assign s_1108 = s_1109 + s_1110;
  assign s_1109 = s_1098?s_1099:s_1101;
  assign s_1110 = s_92 << s_1111;
  assign s_1111 = 5'd29;
  assign s_1112 = 57'd72057594037927936;
  assign s_1113 = 109'd134217728;
  assign s_1114 = s_1115 <= s_155;
  assign s_1115 = s_1116 | s_1120;
  assign s_1116 = s_1117 + s_1118;
  assign s_1117 = s_1106?s_1107:s_1109;
  assign s_1118 = s_90 << s_1119;
  assign s_1119 = 5'd28;
  assign s_1120 = 55'd18014398509481984;
  assign s_1121 = 109'd67108864;
  assign s_1122 = s_1123 <= s_155;
  assign s_1123 = s_1124 | s_1128;
  assign s_1124 = s_1125 + s_1126;
  assign s_1125 = s_1114?s_1115:s_1117;
  assign s_1126 = s_88 << s_1127;
  assign s_1127 = 5'd27;
  assign s_1128 = 53'd4503599627370496;
  assign s_1129 = 109'd33554432;
  assign s_1130 = s_1131 <= s_155;
  assign s_1131 = s_1132 | s_1136;
  assign s_1132 = s_1133 + s_1134;
  assign s_1133 = s_1122?s_1123:s_1125;
  assign s_1134 = s_86 << s_1135;
  assign s_1135 = 5'd26;
  assign s_1136 = 51'd1125899906842624;
  assign s_1137 = 109'd16777216;
  assign s_1138 = s_1139 <= s_155;
  assign s_1139 = s_1140 | s_1144;
  assign s_1140 = s_1141 + s_1142;
  assign s_1141 = s_1130?s_1131:s_1133;
  assign s_1142 = s_84 << s_1143;
  assign s_1143 = 5'd25;
  assign s_1144 = 49'd281474976710656;
  assign s_1145 = 109'd8388608;
  assign s_1146 = s_1147 <= s_155;
  assign s_1147 = s_1148 | s_1152;
  assign s_1148 = s_1149 + s_1150;
  assign s_1149 = s_1138?s_1139:s_1141;
  assign s_1150 = s_82 << s_1151;
  assign s_1151 = 5'd24;
  assign s_1152 = 47'd70368744177664;
  assign s_1153 = 109'd4194304;
  assign s_1154 = s_1155 <= s_155;
  assign s_1155 = s_1156 | s_1160;
  assign s_1156 = s_1157 + s_1158;
  assign s_1157 = s_1146?s_1147:s_1149;
  assign s_1158 = s_80 << s_1159;
  assign s_1159 = 5'd23;
  assign s_1160 = 45'd17592186044416;
  assign s_1161 = 109'd2097152;
  assign s_1162 = s_1163 <= s_155;
  assign s_1163 = s_1164 | s_1168;
  assign s_1164 = s_1165 + s_1166;
  assign s_1165 = s_1154?s_1155:s_1157;
  assign s_1166 = s_78 << s_1167;
  assign s_1167 = 5'd22;
  assign s_1168 = 43'd4398046511104;
  assign s_1169 = 109'd1048576;
  assign s_1170 = s_1171 <= s_155;
  assign s_1171 = s_1172 | s_1176;
  assign s_1172 = s_1173 + s_1174;
  assign s_1173 = s_1162?s_1163:s_1165;
  assign s_1174 = s_76 << s_1175;
  assign s_1175 = 5'd21;
  assign s_1176 = 41'd1099511627776;
  assign s_1177 = 109'd524288;
  assign s_1178 = s_1179 <= s_155;
  assign s_1179 = s_1180 | s_1184;
  assign s_1180 = s_1181 + s_1182;
  assign s_1181 = s_1170?s_1171:s_1173;
  assign s_1182 = s_74 << s_1183;
  assign s_1183 = 5'd20;
  assign s_1184 = 39'd274877906944;
  assign s_1185 = 109'd262144;
  assign s_1186 = s_1187 <= s_155;
  assign s_1187 = s_1188 | s_1192;
  assign s_1188 = s_1189 + s_1190;
  assign s_1189 = s_1178?s_1179:s_1181;
  assign s_1190 = s_72 << s_1191;
  assign s_1191 = 5'd19;
  assign s_1192 = 37'd68719476736;
  assign s_1193 = 109'd131072;
  assign s_1194 = s_1195 <= s_155;
  assign s_1195 = s_1196 | s_1200;
  assign s_1196 = s_1197 + s_1198;
  assign s_1197 = s_1186?s_1187:s_1189;
  assign s_1198 = s_70 << s_1199;
  assign s_1199 = 5'd18;
  assign s_1200 = 35'd17179869184;
  assign s_1201 = 109'd65536;
  assign s_1202 = s_1203 <= s_155;
  assign s_1203 = s_1204 | s_1208;
  assign s_1204 = s_1205 + s_1206;
  assign s_1205 = s_1194?s_1195:s_1197;
  assign s_1206 = s_68 << s_1207;
  assign s_1207 = 5'd17;
  assign s_1208 = 33'd4294967296;
  assign s_1209 = 109'd32768;
  assign s_1210 = s_1211 <= s_155;
  assign s_1211 = s_1212 | s_1216;
  assign s_1212 = s_1213 + s_1214;
  assign s_1213 = s_1202?s_1203:s_1205;
  assign s_1214 = s_66 << s_1215;
  assign s_1215 = 5'd16;
  assign s_1216 = 31'd1073741824;
  assign s_1217 = 109'd16384;
  assign s_1218 = s_1219 <= s_155;
  assign s_1219 = s_1220 | s_1224;
  assign s_1220 = s_1221 + s_1222;
  assign s_1221 = s_1210?s_1211:s_1213;
  assign s_1222 = s_64 << s_1223;
  assign s_1223 = 4'd15;
  assign s_1224 = 29'd268435456;
  assign s_1225 = 109'd8192;
  assign s_1226 = s_1227 <= s_155;
  assign s_1227 = s_1228 | s_1232;
  assign s_1228 = s_1229 + s_1230;
  assign s_1229 = s_1218?s_1219:s_1221;
  assign s_1230 = s_62 << s_1231;
  assign s_1231 = 4'd14;
  assign s_1232 = 27'd67108864;
  assign s_1233 = 109'd4096;
  assign s_1234 = s_1235 <= s_155;
  assign s_1235 = s_1236 | s_1240;
  assign s_1236 = s_1237 + s_1238;
  assign s_1237 = s_1226?s_1227:s_1229;
  assign s_1238 = s_60 << s_1239;
  assign s_1239 = 4'd13;
  assign s_1240 = 25'd16777216;
  assign s_1241 = 109'd2048;
  assign s_1242 = s_1243 <= s_155;
  assign s_1243 = s_1244 | s_1248;
  assign s_1244 = s_1245 + s_1246;
  assign s_1245 = s_1234?s_1235:s_1237;
  assign s_1246 = s_58 << s_1247;
  assign s_1247 = 4'd12;
  assign s_1248 = 23'd4194304;
  assign s_1249 = 109'd1024;
  assign s_1250 = s_1251 <= s_155;
  assign s_1251 = s_1252 | s_1256;
  assign s_1252 = s_1253 + s_1254;
  assign s_1253 = s_1242?s_1243:s_1245;
  assign s_1254 = s_56 << s_1255;
  assign s_1255 = 4'd11;
  assign s_1256 = 21'd1048576;
  assign s_1257 = 109'd512;
  assign s_1258 = s_1259 <= s_155;
  assign s_1259 = s_1260 | s_1264;
  assign s_1260 = s_1261 + s_1262;
  assign s_1261 = s_1250?s_1251:s_1253;
  assign s_1262 = s_54 << s_1263;
  assign s_1263 = 4'd10;
  assign s_1264 = 19'd262144;
  assign s_1265 = 109'd256;
  assign s_1266 = s_1267 <= s_155;
  assign s_1267 = s_1268 | s_1272;
  assign s_1268 = s_1269 + s_1270;
  assign s_1269 = s_1258?s_1259:s_1261;
  assign s_1270 = s_52 << s_1271;
  assign s_1271 = 4'd9;
  assign s_1272 = 17'd65536;
  assign s_1273 = 109'd128;
  assign s_1274 = s_1275 <= s_155;
  assign s_1275 = s_1276 | s_1280;
  assign s_1276 = s_1277 + s_1278;
  assign s_1277 = s_1266?s_1267:s_1269;
  assign s_1278 = s_50 << s_1279;
  assign s_1279 = 4'd8;
  assign s_1280 = 15'd16384;
  assign s_1281 = 109'd64;
  assign s_1282 = s_1283 <= s_155;
  assign s_1283 = s_1284 | s_1288;
  assign s_1284 = s_1285 + s_1286;
  assign s_1285 = s_1274?s_1275:s_1277;
  assign s_1286 = s_48 << s_1287;
  assign s_1287 = 3'd7;
  assign s_1288 = 13'd4096;
  assign s_1289 = 109'd32;
  assign s_1290 = s_1291 <= s_155;
  assign s_1291 = s_1292 | s_1296;
  assign s_1292 = s_1293 + s_1294;
  assign s_1293 = s_1282?s_1283:s_1285;
  assign s_1294 = s_46 << s_1295;
  assign s_1295 = 3'd6;
  assign s_1296 = 11'd1024;
  assign s_1297 = 109'd16;
  assign s_1298 = s_1299 <= s_155;
  assign s_1299 = s_1300 | s_1304;
  assign s_1300 = s_1301 + s_1302;
  assign s_1301 = s_1290?s_1291:s_1293;
  assign s_1302 = s_44 << s_1303;
  assign s_1303 = 3'd5;
  assign s_1304 = 9'd256;
  assign s_1305 = 109'd8;
  assign s_1306 = s_1307 <= s_155;
  assign s_1307 = s_1308 | s_1312;
  assign s_1308 = s_1309 + s_1310;
  assign s_1309 = s_1298?s_1299:s_1301;
  assign s_1310 = s_42 << s_1311;
  assign s_1311 = 3'd4;
  assign s_1312 = 7'd64;
  assign s_1313 = 109'd4;
  assign s_1314 = s_1315 <= s_155;
  assign s_1315 = s_1316 | s_1320;
  assign s_1316 = s_1317 + s_1318;
  assign s_1317 = s_1306?s_1307:s_1309;
  assign s_1318 = s_40 << s_1319;
  assign s_1319 = 2'd3;
  assign s_1320 = 5'd16;
  assign s_1321 = 109'd2;
  assign s_1322 = s_1323 <= s_155;
  assign s_1323 = s_1324 | s_1328;
  assign s_1324 = s_1325 + s_1326;
  assign s_1325 = s_1314?s_1315:s_1317;
  assign s_1326 = s_38 << s_1327;
  assign s_1327 = 2'd2;
  assign s_1328 = 3'd4;
  assign s_1329 = 109'd1;
  assign s_1330 = s_1331 <= s_155;
  assign s_1331 = s_1332 | s_1336;
  assign s_1332 = s_1333 + s_1334;
  assign s_1333 = s_1322?s_1323:s_1325;
  assign s_1334 = s_36 << s_1335;
  assign s_1335 = 1'd1;
  assign s_1336 = 1'd1;
  dq #(13, 1) dq_s_1337 (clk, s_1337, s_1338);
  assign s_1338 = s_1348?s_1339:s_1340;
  assign s_1339 = 1'd0;
  assign s_1340 = s_1341 - s_1342;
  assign s_1341 = -13'd1022;
  dq #(13, 1) dq_s_1342 (clk, s_1342, s_1343);
  assign s_1343 = $signed(s_1344) >>> $signed(s_1347);
  assign s_1344 = s_899?s_1345:s_900;
  assign s_1345 = s_900 - s_1346;
  assign s_1346 = 1'd1;
  assign s_1347 = 13'd1;
  assign s_1348 = s_1340[12];
  dq #(13, 1) dq_s_1349 (clk, s_1349, s_1350);
  assign s_1350 = s_2070?s_1351:s_2064;
  dq #(7, 1) dq_s_1351 (clk, s_1351, s_1352);
  assign s_1352 = {s_1353,s_2058};
  assign s_1353 = s_1354 & s_1716;
  assign s_1354 = s_1355[5];
  assign s_1355 = {s_1356,s_1710};
  assign s_1356 = s_1357 & s_1544;
  assign s_1357 = s_1358[4];
  assign s_1358 = {s_1359,s_1538};
  assign s_1359 = s_1360 & s_1460;
  assign s_1360 = s_1361[3];
  assign s_1361 = {s_1362,s_1454};
  assign s_1362 = s_1363 & s_1420;
  assign s_1363 = s_1364[2];
  assign s_1364 = {s_1365,s_1414};
  assign s_1365 = s_1366 & s_1402;
  assign s_1366 = s_1367[1];
  assign s_1367 = {s_1368,s_1398};
  assign s_1368 = s_1369 & s_1396;
  assign s_1369 = ~s_1370;
  assign s_1370 = s_1371[1];
  assign s_1371 = s_1372[3:2];
  assign s_1372 = s_1373[7:4];
  assign s_1373 = s_1374[15:8];
  assign s_1374 = s_1375[31:16];
  assign s_1375 = s_1376[63:32];
  assign s_1376 = {s_1377,s_1395};
  assign s_1377 = {s_1378,s_1394};
  assign s_1378 = {s_1379,s_1393};
  assign s_1379 = {s_1380,s_1392};
  assign s_1380 = {s_1381,s_1391};
  assign s_1381 = {s_1382,s_1390};
  assign s_1382 = {s_1383,s_1389};
  assign s_1383 = {s_1384,s_1388};
  assign s_1384 = {s_1385,s_1387};
  assign s_1385 = {s_30,s_1386};
  assign s_1386 = 1'd1;
  assign s_1387 = 1'd1;
  assign s_1388 = 1'd1;
  assign s_1389 = 1'd1;
  assign s_1390 = 1'd1;
  assign s_1391 = 1'd1;
  assign s_1392 = 1'd1;
  assign s_1393 = 1'd1;
  assign s_1394 = 1'd1;
  assign s_1395 = 1'd1;
  assign s_1396 = ~s_1397;
  assign s_1397 = s_1371[0];
  assign s_1398 = s_1399 & s_1401;
  assign s_1399 = ~s_1400;
  assign s_1400 = s_1371[1];
  assign s_1401 = s_1371[0];
  assign s_1402 = s_1403[1];
  assign s_1403 = {s_1404,s_1410};
  assign s_1404 = s_1405 & s_1408;
  assign s_1405 = ~s_1406;
  assign s_1406 = s_1407[1];
  assign s_1407 = s_1372[1:0];
  assign s_1408 = ~s_1409;
  assign s_1409 = s_1407[0];
  assign s_1410 = s_1411 & s_1413;
  assign s_1411 = ~s_1412;
  assign s_1412 = s_1407[1];
  assign s_1413 = s_1407[0];
  assign s_1414 = {s_1415,s_1417};
  assign s_1415 = s_1366 & s_1416;
  assign s_1416 = ~s_1402;
  assign s_1417 = s_1366?s_1418:s_1419;
  assign s_1418 = s_1403[0:0];
  assign s_1419 = s_1367[0:0];
  assign s_1420 = s_1421[2];
  assign s_1421 = {s_1422,s_1448};
  assign s_1422 = s_1423 & s_1436;
  assign s_1423 = s_1424[1];
  assign s_1424 = {s_1425,s_1432};
  assign s_1425 = s_1426 & s_1430;
  assign s_1426 = ~s_1427;
  assign s_1427 = s_1428[1];
  assign s_1428 = s_1429[3:2];
  assign s_1429 = s_1373[3:0];
  assign s_1430 = ~s_1431;
  assign s_1431 = s_1428[0];
  assign s_1432 = s_1433 & s_1435;
  assign s_1433 = ~s_1434;
  assign s_1434 = s_1428[1];
  assign s_1435 = s_1428[0];
  assign s_1436 = s_1437[1];
  assign s_1437 = {s_1438,s_1444};
  assign s_1438 = s_1439 & s_1442;
  assign s_1439 = ~s_1440;
  assign s_1440 = s_1441[1];
  assign s_1441 = s_1429[1:0];
  assign s_1442 = ~s_1443;
  assign s_1443 = s_1441[0];
  assign s_1444 = s_1445 & s_1447;
  assign s_1445 = ~s_1446;
  assign s_1446 = s_1441[1];
  assign s_1447 = s_1441[0];
  assign s_1448 = {s_1449,s_1451};
  assign s_1449 = s_1423 & s_1450;
  assign s_1450 = ~s_1436;
  assign s_1451 = s_1423?s_1452:s_1453;
  assign s_1452 = s_1437[0:0];
  assign s_1453 = s_1424[0:0];
  assign s_1454 = {s_1455,s_1457};
  assign s_1455 = s_1363 & s_1456;
  assign s_1456 = ~s_1420;
  assign s_1457 = s_1363?s_1458:s_1459;
  assign s_1458 = s_1421[1:0];
  assign s_1459 = s_1364[1:0];
  assign s_1460 = s_1461[3];
  assign s_1461 = {s_1462,s_1532};
  assign s_1462 = s_1463 & s_1498;
  assign s_1463 = s_1464[2];
  assign s_1464 = {s_1465,s_1492};
  assign s_1465 = s_1466 & s_1480;
  assign s_1466 = s_1467[1];
  assign s_1467 = {s_1468,s_1476};
  assign s_1468 = s_1469 & s_1474;
  assign s_1469 = ~s_1470;
  assign s_1470 = s_1471[1];
  assign s_1471 = s_1472[3:2];
  assign s_1472 = s_1473[7:4];
  assign s_1473 = s_1374[7:0];
  assign s_1474 = ~s_1475;
  assign s_1475 = s_1471[0];
  assign s_1476 = s_1477 & s_1479;
  assign s_1477 = ~s_1478;
  assign s_1478 = s_1471[1];
  assign s_1479 = s_1471[0];
  assign s_1480 = s_1481[1];
  assign s_1481 = {s_1482,s_1488};
  assign s_1482 = s_1483 & s_1486;
  assign s_1483 = ~s_1484;
  assign s_1484 = s_1485[1];
  assign s_1485 = s_1472[1:0];
  assign s_1486 = ~s_1487;
  assign s_1487 = s_1485[0];
  assign s_1488 = s_1489 & s_1491;
  assign s_1489 = ~s_1490;
  assign s_1490 = s_1485[1];
  assign s_1491 = s_1485[0];
  assign s_1492 = {s_1493,s_1495};
  assign s_1493 = s_1466 & s_1494;
  assign s_1494 = ~s_1480;
  assign s_1495 = s_1466?s_1496:s_1497;
  assign s_1496 = s_1481[0:0];
  assign s_1497 = s_1467[0:0];
  assign s_1498 = s_1499[2];
  assign s_1499 = {s_1500,s_1526};
  assign s_1500 = s_1501 & s_1514;
  assign s_1501 = s_1502[1];
  assign s_1502 = {s_1503,s_1510};
  assign s_1503 = s_1504 & s_1508;
  assign s_1504 = ~s_1505;
  assign s_1505 = s_1506[1];
  assign s_1506 = s_1507[3:2];
  assign s_1507 = s_1473[3:0];
  assign s_1508 = ~s_1509;
  assign s_1509 = s_1506[0];
  assign s_1510 = s_1511 & s_1513;
  assign s_1511 = ~s_1512;
  assign s_1512 = s_1506[1];
  assign s_1513 = s_1506[0];
  assign s_1514 = s_1515[1];
  assign s_1515 = {s_1516,s_1522};
  assign s_1516 = s_1517 & s_1520;
  assign s_1517 = ~s_1518;
  assign s_1518 = s_1519[1];
  assign s_1519 = s_1507[1:0];
  assign s_1520 = ~s_1521;
  assign s_1521 = s_1519[0];
  assign s_1522 = s_1523 & s_1525;
  assign s_1523 = ~s_1524;
  assign s_1524 = s_1519[1];
  assign s_1525 = s_1519[0];
  assign s_1526 = {s_1527,s_1529};
  assign s_1527 = s_1501 & s_1528;
  assign s_1528 = ~s_1514;
  assign s_1529 = s_1501?s_1530:s_1531;
  assign s_1530 = s_1515[0:0];
  assign s_1531 = s_1502[0:0];
  assign s_1532 = {s_1533,s_1535};
  assign s_1533 = s_1463 & s_1534;
  assign s_1534 = ~s_1498;
  assign s_1535 = s_1463?s_1536:s_1537;
  assign s_1536 = s_1499[1:0];
  assign s_1537 = s_1464[1:0];
  assign s_1538 = {s_1539,s_1541};
  assign s_1539 = s_1360 & s_1540;
  assign s_1540 = ~s_1460;
  assign s_1541 = s_1360?s_1542:s_1543;
  assign s_1542 = s_1461[2:0];
  assign s_1543 = s_1361[2:0];
  assign s_1544 = s_1545[4];
  assign s_1545 = {s_1546,s_1704};
  assign s_1546 = s_1547 & s_1626;
  assign s_1547 = s_1548[3];
  assign s_1548 = {s_1549,s_1620};
  assign s_1549 = s_1550 & s_1586;
  assign s_1550 = s_1551[2];
  assign s_1551 = {s_1552,s_1580};
  assign s_1552 = s_1553 & s_1568;
  assign s_1553 = s_1554[1];
  assign s_1554 = {s_1555,s_1564};
  assign s_1555 = s_1556 & s_1562;
  assign s_1556 = ~s_1557;
  assign s_1557 = s_1558[1];
  assign s_1558 = s_1559[3:2];
  assign s_1559 = s_1560[7:4];
  assign s_1560 = s_1561[15:8];
  assign s_1561 = s_1375[15:0];
  assign s_1562 = ~s_1563;
  assign s_1563 = s_1558[0];
  assign s_1564 = s_1565 & s_1567;
  assign s_1565 = ~s_1566;
  assign s_1566 = s_1558[1];
  assign s_1567 = s_1558[0];
  assign s_1568 = s_1569[1];
  assign s_1569 = {s_1570,s_1576};
  assign s_1570 = s_1571 & s_1574;
  assign s_1571 = ~s_1572;
  assign s_1572 = s_1573[1];
  assign s_1573 = s_1559[1:0];
  assign s_1574 = ~s_1575;
  assign s_1575 = s_1573[0];
  assign s_1576 = s_1577 & s_1579;
  assign s_1577 = ~s_1578;
  assign s_1578 = s_1573[1];
  assign s_1579 = s_1573[0];
  assign s_1580 = {s_1581,s_1583};
  assign s_1581 = s_1553 & s_1582;
  assign s_1582 = ~s_1568;
  assign s_1583 = s_1553?s_1584:s_1585;
  assign s_1584 = s_1569[0:0];
  assign s_1585 = s_1554[0:0];
  assign s_1586 = s_1587[2];
  assign s_1587 = {s_1588,s_1614};
  assign s_1588 = s_1589 & s_1602;
  assign s_1589 = s_1590[1];
  assign s_1590 = {s_1591,s_1598};
  assign s_1591 = s_1592 & s_1596;
  assign s_1592 = ~s_1593;
  assign s_1593 = s_1594[1];
  assign s_1594 = s_1595[3:2];
  assign s_1595 = s_1560[3:0];
  assign s_1596 = ~s_1597;
  assign s_1597 = s_1594[0];
  assign s_1598 = s_1599 & s_1601;
  assign s_1599 = ~s_1600;
  assign s_1600 = s_1594[1];
  assign s_1601 = s_1594[0];
  assign s_1602 = s_1603[1];
  assign s_1603 = {s_1604,s_1610};
  assign s_1604 = s_1605 & s_1608;
  assign s_1605 = ~s_1606;
  assign s_1606 = s_1607[1];
  assign s_1607 = s_1595[1:0];
  assign s_1608 = ~s_1609;
  assign s_1609 = s_1607[0];
  assign s_1610 = s_1611 & s_1613;
  assign s_1611 = ~s_1612;
  assign s_1612 = s_1607[1];
  assign s_1613 = s_1607[0];
  assign s_1614 = {s_1615,s_1617};
  assign s_1615 = s_1589 & s_1616;
  assign s_1616 = ~s_1602;
  assign s_1617 = s_1589?s_1618:s_1619;
  assign s_1618 = s_1603[0:0];
  assign s_1619 = s_1590[0:0];
  assign s_1620 = {s_1621,s_1623};
  assign s_1621 = s_1550 & s_1622;
  assign s_1622 = ~s_1586;
  assign s_1623 = s_1550?s_1624:s_1625;
  assign s_1624 = s_1587[1:0];
  assign s_1625 = s_1551[1:0];
  assign s_1626 = s_1627[3];
  assign s_1627 = {s_1628,s_1698};
  assign s_1628 = s_1629 & s_1664;
  assign s_1629 = s_1630[2];
  assign s_1630 = {s_1631,s_1658};
  assign s_1631 = s_1632 & s_1646;
  assign s_1632 = s_1633[1];
  assign s_1633 = {s_1634,s_1642};
  assign s_1634 = s_1635 & s_1640;
  assign s_1635 = ~s_1636;
  assign s_1636 = s_1637[1];
  assign s_1637 = s_1638[3:2];
  assign s_1638 = s_1639[7:4];
  assign s_1639 = s_1561[7:0];
  assign s_1640 = ~s_1641;
  assign s_1641 = s_1637[0];
  assign s_1642 = s_1643 & s_1645;
  assign s_1643 = ~s_1644;
  assign s_1644 = s_1637[1];
  assign s_1645 = s_1637[0];
  assign s_1646 = s_1647[1];
  assign s_1647 = {s_1648,s_1654};
  assign s_1648 = s_1649 & s_1652;
  assign s_1649 = ~s_1650;
  assign s_1650 = s_1651[1];
  assign s_1651 = s_1638[1:0];
  assign s_1652 = ~s_1653;
  assign s_1653 = s_1651[0];
  assign s_1654 = s_1655 & s_1657;
  assign s_1655 = ~s_1656;
  assign s_1656 = s_1651[1];
  assign s_1657 = s_1651[0];
  assign s_1658 = {s_1659,s_1661};
  assign s_1659 = s_1632 & s_1660;
  assign s_1660 = ~s_1646;
  assign s_1661 = s_1632?s_1662:s_1663;
  assign s_1662 = s_1647[0:0];
  assign s_1663 = s_1633[0:0];
  assign s_1664 = s_1665[2];
  assign s_1665 = {s_1666,s_1692};
  assign s_1666 = s_1667 & s_1680;
  assign s_1667 = s_1668[1];
  assign s_1668 = {s_1669,s_1676};
  assign s_1669 = s_1670 & s_1674;
  assign s_1670 = ~s_1671;
  assign s_1671 = s_1672[1];
  assign s_1672 = s_1673[3:2];
  assign s_1673 = s_1639[3:0];
  assign s_1674 = ~s_1675;
  assign s_1675 = s_1672[0];
  assign s_1676 = s_1677 & s_1679;
  assign s_1677 = ~s_1678;
  assign s_1678 = s_1672[1];
  assign s_1679 = s_1672[0];
  assign s_1680 = s_1681[1];
  assign s_1681 = {s_1682,s_1688};
  assign s_1682 = s_1683 & s_1686;
  assign s_1683 = ~s_1684;
  assign s_1684 = s_1685[1];
  assign s_1685 = s_1673[1:0];
  assign s_1686 = ~s_1687;
  assign s_1687 = s_1685[0];
  assign s_1688 = s_1689 & s_1691;
  assign s_1689 = ~s_1690;
  assign s_1690 = s_1685[1];
  assign s_1691 = s_1685[0];
  assign s_1692 = {s_1693,s_1695};
  assign s_1693 = s_1667 & s_1694;
  assign s_1694 = ~s_1680;
  assign s_1695 = s_1667?s_1696:s_1697;
  assign s_1696 = s_1681[0:0];
  assign s_1697 = s_1668[0:0];
  assign s_1698 = {s_1699,s_1701};
  assign s_1699 = s_1629 & s_1700;
  assign s_1700 = ~s_1664;
  assign s_1701 = s_1629?s_1702:s_1703;
  assign s_1702 = s_1665[1:0];
  assign s_1703 = s_1630[1:0];
  assign s_1704 = {s_1705,s_1707};
  assign s_1705 = s_1547 & s_1706;
  assign s_1706 = ~s_1626;
  assign s_1707 = s_1547?s_1708:s_1709;
  assign s_1708 = s_1627[2:0];
  assign s_1709 = s_1548[2:0];
  assign s_1710 = {s_1711,s_1713};
  assign s_1711 = s_1357 & s_1712;
  assign s_1712 = ~s_1544;
  assign s_1713 = s_1357?s_1714:s_1715;
  assign s_1714 = s_1545[3:0];
  assign s_1715 = s_1358[3:0];
  assign s_1716 = s_1717[5];
  assign s_1717 = {s_1718,s_2052};
  assign s_1718 = s_1719 & s_1886;
  assign s_1719 = s_1720[4];
  assign s_1720 = {s_1721,s_1880};
  assign s_1721 = s_1722 & s_1802;
  assign s_1722 = s_1723[3];
  assign s_1723 = {s_1724,s_1796};
  assign s_1724 = s_1725 & s_1762;
  assign s_1725 = s_1726[2];
  assign s_1726 = {s_1727,s_1756};
  assign s_1727 = s_1728 & s_1744;
  assign s_1728 = s_1729[1];
  assign s_1729 = {s_1730,s_1740};
  assign s_1730 = s_1731 & s_1738;
  assign s_1731 = ~s_1732;
  assign s_1732 = s_1733[1];
  assign s_1733 = s_1734[3:2];
  assign s_1734 = s_1735[7:4];
  assign s_1735 = s_1736[15:8];
  assign s_1736 = s_1737[31:16];
  assign s_1737 = s_1376[31:0];
  assign s_1738 = ~s_1739;
  assign s_1739 = s_1733[0];
  assign s_1740 = s_1741 & s_1743;
  assign s_1741 = ~s_1742;
  assign s_1742 = s_1733[1];
  assign s_1743 = s_1733[0];
  assign s_1744 = s_1745[1];
  assign s_1745 = {s_1746,s_1752};
  assign s_1746 = s_1747 & s_1750;
  assign s_1747 = ~s_1748;
  assign s_1748 = s_1749[1];
  assign s_1749 = s_1734[1:0];
  assign s_1750 = ~s_1751;
  assign s_1751 = s_1749[0];
  assign s_1752 = s_1753 & s_1755;
  assign s_1753 = ~s_1754;
  assign s_1754 = s_1749[1];
  assign s_1755 = s_1749[0];
  assign s_1756 = {s_1757,s_1759};
  assign s_1757 = s_1728 & s_1758;
  assign s_1758 = ~s_1744;
  assign s_1759 = s_1728?s_1760:s_1761;
  assign s_1760 = s_1745[0:0];
  assign s_1761 = s_1729[0:0];
  assign s_1762 = s_1763[2];
  assign s_1763 = {s_1764,s_1790};
  assign s_1764 = s_1765 & s_1778;
  assign s_1765 = s_1766[1];
  assign s_1766 = {s_1767,s_1774};
  assign s_1767 = s_1768 & s_1772;
  assign s_1768 = ~s_1769;
  assign s_1769 = s_1770[1];
  assign s_1770 = s_1771[3:2];
  assign s_1771 = s_1735[3:0];
  assign s_1772 = ~s_1773;
  assign s_1773 = s_1770[0];
  assign s_1774 = s_1775 & s_1777;
  assign s_1775 = ~s_1776;
  assign s_1776 = s_1770[1];
  assign s_1777 = s_1770[0];
  assign s_1778 = s_1779[1];
  assign s_1779 = {s_1780,s_1786};
  assign s_1780 = s_1781 & s_1784;
  assign s_1781 = ~s_1782;
  assign s_1782 = s_1783[1];
  assign s_1783 = s_1771[1:0];
  assign s_1784 = ~s_1785;
  assign s_1785 = s_1783[0];
  assign s_1786 = s_1787 & s_1789;
  assign s_1787 = ~s_1788;
  assign s_1788 = s_1783[1];
  assign s_1789 = s_1783[0];
  assign s_1790 = {s_1791,s_1793};
  assign s_1791 = s_1765 & s_1792;
  assign s_1792 = ~s_1778;
  assign s_1793 = s_1765?s_1794:s_1795;
  assign s_1794 = s_1779[0:0];
  assign s_1795 = s_1766[0:0];
  assign s_1796 = {s_1797,s_1799};
  assign s_1797 = s_1725 & s_1798;
  assign s_1798 = ~s_1762;
  assign s_1799 = s_1725?s_1800:s_1801;
  assign s_1800 = s_1763[1:0];
  assign s_1801 = s_1726[1:0];
  assign s_1802 = s_1803[3];
  assign s_1803 = {s_1804,s_1874};
  assign s_1804 = s_1805 & s_1840;
  assign s_1805 = s_1806[2];
  assign s_1806 = {s_1807,s_1834};
  assign s_1807 = s_1808 & s_1822;
  assign s_1808 = s_1809[1];
  assign s_1809 = {s_1810,s_1818};
  assign s_1810 = s_1811 & s_1816;
  assign s_1811 = ~s_1812;
  assign s_1812 = s_1813[1];
  assign s_1813 = s_1814[3:2];
  assign s_1814 = s_1815[7:4];
  assign s_1815 = s_1736[7:0];
  assign s_1816 = ~s_1817;
  assign s_1817 = s_1813[0];
  assign s_1818 = s_1819 & s_1821;
  assign s_1819 = ~s_1820;
  assign s_1820 = s_1813[1];
  assign s_1821 = s_1813[0];
  assign s_1822 = s_1823[1];
  assign s_1823 = {s_1824,s_1830};
  assign s_1824 = s_1825 & s_1828;
  assign s_1825 = ~s_1826;
  assign s_1826 = s_1827[1];
  assign s_1827 = s_1814[1:0];
  assign s_1828 = ~s_1829;
  assign s_1829 = s_1827[0];
  assign s_1830 = s_1831 & s_1833;
  assign s_1831 = ~s_1832;
  assign s_1832 = s_1827[1];
  assign s_1833 = s_1827[0];
  assign s_1834 = {s_1835,s_1837};
  assign s_1835 = s_1808 & s_1836;
  assign s_1836 = ~s_1822;
  assign s_1837 = s_1808?s_1838:s_1839;
  assign s_1838 = s_1823[0:0];
  assign s_1839 = s_1809[0:0];
  assign s_1840 = s_1841[2];
  assign s_1841 = {s_1842,s_1868};
  assign s_1842 = s_1843 & s_1856;
  assign s_1843 = s_1844[1];
  assign s_1844 = {s_1845,s_1852};
  assign s_1845 = s_1846 & s_1850;
  assign s_1846 = ~s_1847;
  assign s_1847 = s_1848[1];
  assign s_1848 = s_1849[3:2];
  assign s_1849 = s_1815[3:0];
  assign s_1850 = ~s_1851;
  assign s_1851 = s_1848[0];
  assign s_1852 = s_1853 & s_1855;
  assign s_1853 = ~s_1854;
  assign s_1854 = s_1848[1];
  assign s_1855 = s_1848[0];
  assign s_1856 = s_1857[1];
  assign s_1857 = {s_1858,s_1864};
  assign s_1858 = s_1859 & s_1862;
  assign s_1859 = ~s_1860;
  assign s_1860 = s_1861[1];
  assign s_1861 = s_1849[1:0];
  assign s_1862 = ~s_1863;
  assign s_1863 = s_1861[0];
  assign s_1864 = s_1865 & s_1867;
  assign s_1865 = ~s_1866;
  assign s_1866 = s_1861[1];
  assign s_1867 = s_1861[0];
  assign s_1868 = {s_1869,s_1871};
  assign s_1869 = s_1843 & s_1870;
  assign s_1870 = ~s_1856;
  assign s_1871 = s_1843?s_1872:s_1873;
  assign s_1872 = s_1857[0:0];
  assign s_1873 = s_1844[0:0];
  assign s_1874 = {s_1875,s_1877};
  assign s_1875 = s_1805 & s_1876;
  assign s_1876 = ~s_1840;
  assign s_1877 = s_1805?s_1878:s_1879;
  assign s_1878 = s_1841[1:0];
  assign s_1879 = s_1806[1:0];
  assign s_1880 = {s_1881,s_1883};
  assign s_1881 = s_1722 & s_1882;
  assign s_1882 = ~s_1802;
  assign s_1883 = s_1722?s_1884:s_1885;
  assign s_1884 = s_1803[2:0];
  assign s_1885 = s_1723[2:0];
  assign s_1886 = s_1887[4];
  assign s_1887 = {s_1888,s_2046};
  assign s_1888 = s_1889 & s_1968;
  assign s_1889 = s_1890[3];
  assign s_1890 = {s_1891,s_1962};
  assign s_1891 = s_1892 & s_1928;
  assign s_1892 = s_1893[2];
  assign s_1893 = {s_1894,s_1922};
  assign s_1894 = s_1895 & s_1910;
  assign s_1895 = s_1896[1];
  assign s_1896 = {s_1897,s_1906};
  assign s_1897 = s_1898 & s_1904;
  assign s_1898 = ~s_1899;
  assign s_1899 = s_1900[1];
  assign s_1900 = s_1901[3:2];
  assign s_1901 = s_1902[7:4];
  assign s_1902 = s_1903[15:8];
  assign s_1903 = s_1737[15:0];
  assign s_1904 = ~s_1905;
  assign s_1905 = s_1900[0];
  assign s_1906 = s_1907 & s_1909;
  assign s_1907 = ~s_1908;
  assign s_1908 = s_1900[1];
  assign s_1909 = s_1900[0];
  assign s_1910 = s_1911[1];
  assign s_1911 = {s_1912,s_1918};
  assign s_1912 = s_1913 & s_1916;
  assign s_1913 = ~s_1914;
  assign s_1914 = s_1915[1];
  assign s_1915 = s_1901[1:0];
  assign s_1916 = ~s_1917;
  assign s_1917 = s_1915[0];
  assign s_1918 = s_1919 & s_1921;
  assign s_1919 = ~s_1920;
  assign s_1920 = s_1915[1];
  assign s_1921 = s_1915[0];
  assign s_1922 = {s_1923,s_1925};
  assign s_1923 = s_1895 & s_1924;
  assign s_1924 = ~s_1910;
  assign s_1925 = s_1895?s_1926:s_1927;
  assign s_1926 = s_1911[0:0];
  assign s_1927 = s_1896[0:0];
  assign s_1928 = s_1929[2];
  assign s_1929 = {s_1930,s_1956};
  assign s_1930 = s_1931 & s_1944;
  assign s_1931 = s_1932[1];
  assign s_1932 = {s_1933,s_1940};
  assign s_1933 = s_1934 & s_1938;
  assign s_1934 = ~s_1935;
  assign s_1935 = s_1936[1];
  assign s_1936 = s_1937[3:2];
  assign s_1937 = s_1902[3:0];
  assign s_1938 = ~s_1939;
  assign s_1939 = s_1936[0];
  assign s_1940 = s_1941 & s_1943;
  assign s_1941 = ~s_1942;
  assign s_1942 = s_1936[1];
  assign s_1943 = s_1936[0];
  assign s_1944 = s_1945[1];
  assign s_1945 = {s_1946,s_1952};
  assign s_1946 = s_1947 & s_1950;
  assign s_1947 = ~s_1948;
  assign s_1948 = s_1949[1];
  assign s_1949 = s_1937[1:0];
  assign s_1950 = ~s_1951;
  assign s_1951 = s_1949[0];
  assign s_1952 = s_1953 & s_1955;
  assign s_1953 = ~s_1954;
  assign s_1954 = s_1949[1];
  assign s_1955 = s_1949[0];
  assign s_1956 = {s_1957,s_1959};
  assign s_1957 = s_1931 & s_1958;
  assign s_1958 = ~s_1944;
  assign s_1959 = s_1931?s_1960:s_1961;
  assign s_1960 = s_1945[0:0];
  assign s_1961 = s_1932[0:0];
  assign s_1962 = {s_1963,s_1965};
  assign s_1963 = s_1892 & s_1964;
  assign s_1964 = ~s_1928;
  assign s_1965 = s_1892?s_1966:s_1967;
  assign s_1966 = s_1929[1:0];
  assign s_1967 = s_1893[1:0];
  assign s_1968 = s_1969[3];
  assign s_1969 = {s_1970,s_2040};
  assign s_1970 = s_1971 & s_2006;
  assign s_1971 = s_1972[2];
  assign s_1972 = {s_1973,s_2000};
  assign s_1973 = s_1974 & s_1988;
  assign s_1974 = s_1975[1];
  assign s_1975 = {s_1976,s_1984};
  assign s_1976 = s_1977 & s_1982;
  assign s_1977 = ~s_1978;
  assign s_1978 = s_1979[1];
  assign s_1979 = s_1980[3:2];
  assign s_1980 = s_1981[7:4];
  assign s_1981 = s_1903[7:0];
  assign s_1982 = ~s_1983;
  assign s_1983 = s_1979[0];
  assign s_1984 = s_1985 & s_1987;
  assign s_1985 = ~s_1986;
  assign s_1986 = s_1979[1];
  assign s_1987 = s_1979[0];
  assign s_1988 = s_1989[1];
  assign s_1989 = {s_1990,s_1996};
  assign s_1990 = s_1991 & s_1994;
  assign s_1991 = ~s_1992;
  assign s_1992 = s_1993[1];
  assign s_1993 = s_1980[1:0];
  assign s_1994 = ~s_1995;
  assign s_1995 = s_1993[0];
  assign s_1996 = s_1997 & s_1999;
  assign s_1997 = ~s_1998;
  assign s_1998 = s_1993[1];
  assign s_1999 = s_1993[0];
  assign s_2000 = {s_2001,s_2003};
  assign s_2001 = s_1974 & s_2002;
  assign s_2002 = ~s_1988;
  assign s_2003 = s_1974?s_2004:s_2005;
  assign s_2004 = s_1989[0:0];
  assign s_2005 = s_1975[0:0];
  assign s_2006 = s_2007[2];
  assign s_2007 = {s_2008,s_2034};
  assign s_2008 = s_2009 & s_2022;
  assign s_2009 = s_2010[1];
  assign s_2010 = {s_2011,s_2018};
  assign s_2011 = s_2012 & s_2016;
  assign s_2012 = ~s_2013;
  assign s_2013 = s_2014[1];
  assign s_2014 = s_2015[3:2];
  assign s_2015 = s_1981[3:0];
  assign s_2016 = ~s_2017;
  assign s_2017 = s_2014[0];
  assign s_2018 = s_2019 & s_2021;
  assign s_2019 = ~s_2020;
  assign s_2020 = s_2014[1];
  assign s_2021 = s_2014[0];
  assign s_2022 = s_2023[1];
  assign s_2023 = {s_2024,s_2030};
  assign s_2024 = s_2025 & s_2028;
  assign s_2025 = ~s_2026;
  assign s_2026 = s_2027[1];
  assign s_2027 = s_2015[1:0];
  assign s_2028 = ~s_2029;
  assign s_2029 = s_2027[0];
  assign s_2030 = s_2031 & s_2033;
  assign s_2031 = ~s_2032;
  assign s_2032 = s_2027[1];
  assign s_2033 = s_2027[0];
  assign s_2034 = {s_2035,s_2037};
  assign s_2035 = s_2009 & s_2036;
  assign s_2036 = ~s_2022;
  assign s_2037 = s_2009?s_2038:s_2039;
  assign s_2038 = s_2023[0:0];
  assign s_2039 = s_2010[0:0];
  assign s_2040 = {s_2041,s_2043};
  assign s_2041 = s_1971 & s_2042;
  assign s_2042 = ~s_2006;
  assign s_2043 = s_1971?s_2044:s_2045;
  assign s_2044 = s_2007[1:0];
  assign s_2045 = s_1972[1:0];
  assign s_2046 = {s_2047,s_2049};
  assign s_2047 = s_1889 & s_2048;
  assign s_2048 = ~s_1968;
  assign s_2049 = s_1889?s_2050:s_2051;
  assign s_2050 = s_1969[2:0];
  assign s_2051 = s_1890[2:0];
  assign s_2052 = {s_2053,s_2055};
  assign s_2053 = s_1719 & s_2054;
  assign s_2054 = ~s_1886;
  assign s_2055 = s_1719?s_2056:s_2057;
  assign s_2056 = s_1887[3:0];
  assign s_2057 = s_1720[3:0];
  assign s_2058 = {s_2059,s_2061};
  assign s_2059 = s_1354 & s_2060;
  assign s_2060 = ~s_1716;
  assign s_2061 = s_1354?s_2062:s_2063;
  assign s_2062 = s_1717[4:0];
  assign s_2063 = s_1355[4:0];
  dq #(13, 1) dq_s_2064 (clk, s_2064, s_2065);
  assign s_2065 = s_2066 - s_2069;
  dq #(13, 1) dq_s_2066 (clk, s_2066, s_2067);
  assign s_2067 = s_2068 + s_1337;
  dq #(13, 1) dq_s_2068 (clk, s_2068, s_1342);
  assign s_2069 = -13'd1022;
  assign s_2070 = s_2071 <= s_2072;
  assign s_2071 = s_1351;
  dq #(13, 1) dq_s_2072 (clk, s_2072, s_2065);
  assign s_2073 = 1'd1;
  assign s_2074 = s_2075 & s_2076;
  assign s_2075 = s_27[0];
  assign s_2076 = s_2077 | s_2081;
  dq #(1, 9) dq_s_2077 (clk, s_2077, s_2078);
  assign s_2078 = s_2079 | s_2080;
  assign s_2079 = 1'd1;
  assign s_2080 = 1'd0;
  assign s_2081 = s_26[0];
  assign s_2082 = s_23[52:0];
  assign s_2083 = s_23[53];
  assign s_2084 = {s_2085,s_2095};
  assign s_2085 = {s_2086,s_2087};
  dq #(1, 10) dq_s_2086 (clk, s_2086, s_3);
  assign s_2087 = s_2088 + s_2094;
  assign s_2088 = s_2089[10:0];
  dq #(13, 1) dq_s_2089 (clk, s_2089, s_2090);
  assign s_2090 = s_2091 + s_2083;
  dq #(13, 1) dq_s_2091 (clk, s_2091, s_2092);
  assign s_2092 = s_2093 - s_1349;
  dq #(13, 2) dq_s_2093 (clk, s_2093, s_2066);
  assign s_2094 = 10'd1023;
  assign s_2095 = s_20[51:0];
  assign s_2096 = s_2097 & s_2099;
  assign s_2097 = s_2088 == s_2098;
  assign s_2098 = -11'd1022;
  assign s_2099 = ~s_2100;
  assign s_2100 = s_20[52];
  assign s_2101 = s_20 == s_2102;
  assign s_2102 = 53'd0;
  dq #(1, 10) dq_s_2103 (clk, s_2103, s_2104);
  assign s_2104 = s_2105 & s_2107;
  assign s_2105 = s_167 == s_2106;
  assign s_2106 = 11'd1024;
  assign s_2107 = s_171 == s_2108;
  assign s_2108 = 52'd0;
  assign s_2109 = s_2110 | s_2116;
  dq #(1, 10) dq_s_2110 (clk, s_2110, s_2111);
  assign s_2111 = s_2112 & s_2114;
  assign s_2112 = s_167 == s_2113;
  assign s_2113 = 11'd1024;
  assign s_2114 = s_171 != s_2115;
  assign s_2115 = 52'd0;
  assign s_2116 = s_2117 & s_2118;
  dq #(1, 10) dq_s_2117 (clk, s_2117, s_3);
  assign s_2118 = s_20 != s_2119;
  assign s_2119 = 1'd0;
  assign double_sqrt_z = s_0;
endmodule
